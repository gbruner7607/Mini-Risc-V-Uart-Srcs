
// Netlisted models

// Library - sram_compiled_r128_c128_w8, Cell - colDecoder, View -
//schematic
// LAST TIME SAVED: Apr 20 20:07:34 2021
// NETLIST TIME: Apr 21 18:57:09 2021
`timescale 1ns / 1ps 

module colDecoder ( A0, A0_inv, A1, A1_inv, A2, A2_inv, A3, A3_inv,
     CLK, YF0, YF1, YF2, YF3, YF4, YF5, YF6, YF7, YF8, YF9, YF10, YF11,
     YF12, YF13, YF14, YF15 );

output  YF0, YF1, YF2, YF3, YF4, YF5, YF6, YF7, YF8, YF9, YF10, YF11,
     YF12, YF13, YF14, YF15;

input  A0, A0_inv, A1, A1_inv, A2, A2_inv, A3, A3_inv, CLK;


specify 
    specparam CDS_LIBNAME  = "sram_compiled_r128_c128_w8";
    specparam CDS_CELLNAME = "colDecoder";
    specparam CDS_VIEWNAME = "schematic";
endspecify

NANDC2x1 inst_clockedAND_b15_15 ( imd_YF15, CLK, Y15);
NANDC2x1 inst_and_b15_0_1 ( imd_wire15_0_1, A2, A3);
NANDC2x1 inst_and_b15_0_0 ( imd_wire15_0_0, A0, A1);
NANDC2x1 inst_and_b15_1_0 ( imd_Y15, wire15_0_0, wire15_0_1);
NANDC2x1 inst_clockedAND_b14_14 ( imd_YF14, CLK, Y14);
NANDC2x1 inst_and_b14_0_1 ( imd_wire14_0_1, A2, A3);
NANDC2x1 inst_and_b14_0_0 ( imd_wire14_0_0, A0_inv, A1);
NANDC2x1 inst_and_b14_1_0 ( imd_Y14, wire14_0_0, wire14_0_1);
NANDC2x1 inst_clockedAND_b13_13 ( imd_YF13, CLK, Y13);
NANDC2x1 inst_and_b13_0_1 ( imd_wire13_0_1, A2, A3);
NANDC2x1 inst_and_b13_0_0 ( imd_wire13_0_0, A0, A1_inv);
NANDC2x1 inst_and_b13_1_0 ( imd_Y13, wire13_0_0, wire13_0_1);
NANDC2x1 inst_clockedAND_b12_12 ( imd_YF12, CLK, Y12);
NANDC2x1 inst_and_b12_0_1 ( imd_wire12_0_1, A2, A3);
NANDC2x1 inst_and_b12_0_0 ( imd_wire12_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b12_1_0 ( imd_Y12, wire12_0_0, wire12_0_1);
NANDC2x1 inst_clockedAND_b11_11 ( imd_YF11, CLK, Y11);
NANDC2x1 inst_and_b11_0_1 ( imd_wire11_0_1, A2_inv, A3);
NANDC2x1 inst_and_b11_0_0 ( imd_wire11_0_0, A0, A1);
NANDC2x1 inst_and_b11_1_0 ( imd_Y11, wire11_0_0, wire11_0_1);
NANDC2x1 inst_clockedAND_b10_10 ( imd_YF10, CLK, Y10);
NANDC2x1 inst_and_b10_0_1 ( imd_wire10_0_1, A2_inv, A3);
NANDC2x1 inst_and_b10_0_0 ( imd_wire10_0_0, A0_inv, A1);
NANDC2x1 inst_and_b10_1_0 ( imd_Y10, wire10_0_0, wire10_0_1);
NANDC2x1 inst_clockedAND_b9_9 ( imd_YF9, CLK, Y9);
NANDC2x1 inst_and_b9_0_1 ( imd_wire9_0_1, A2_inv, A3);
NANDC2x1 inst_and_b9_0_0 ( imd_wire9_0_0, A0, A1_inv);
NANDC2x1 inst_and_b9_1_0 ( imd_Y9, wire9_0_0, wire9_0_1);
NANDC2x1 inst_and_b8_0_1 ( imd_wire8_0_1, A2_inv, A3);
NANDC2x1 inst_clockedAND_b8_8 ( imd_YF8, CLK, Y8);
NANDC2x1 inst_and_b8_0_0 ( imd_wire8_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b8_1_0 ( imd_Y8, wire8_0_0, wire8_0_1);
NANDC2x1 inst_clockedAND_b7_7 ( imd_YF7, CLK, Y7);
NANDC2x1 inst_and_b7_0_1 ( imd_wire7_0_1, A2, A3_inv);
NANDC2x1 inst_and_b7_0_0 ( imd_wire7_0_0, A0, A1);
NANDC2x1 inst_and_b7_1_0 ( imd_Y7, wire7_0_0, wire7_0_1);
NANDC2x1 inst_clockedAND_b6_6 ( imd_YF6, CLK, Y6);
NANDC2x1 inst_and_b6_0_1 ( imd_wire6_0_1, A2, A3_inv);
NANDC2x1 inst_and_b6_0_0 ( imd_wire6_0_0, A0_inv, A1);
NANDC2x1 inst_and_b6_1_0 ( imd_Y6, wire6_0_0, wire6_0_1);
NANDC2x1 inst_clockedAND_b5_5 ( imd_YF5, CLK, Y5);
NANDC2x1 inst_and_b5_0_1 ( imd_wire5_0_1, A2, A3_inv);
NANDC2x1 inst_and_b5_0_0 ( imd_wire5_0_0, A0, A1_inv);
NANDC2x1 inst_and_b5_1_0 ( imd_Y5, wire5_0_0, wire5_0_1);
NANDC2x1 inst_and_b4_0_1 ( imd_wire4_0_1, A2, A3_inv);
NANDC2x1 inst_clockedAND_b4_4 ( imd_YF4, CLK, Y4);
NANDC2x1 inst_and_b4_0_0 ( imd_wire4_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b4_1_0 ( imd_Y4, wire4_0_0, wire4_0_1);
NANDC2x1 inst_clockedAND_b3_3 ( imd_YF3, CLK, Y3);
NANDC2x1 inst_and_b3_0_1 ( imd_wire3_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b3_0_0 ( imd_wire3_0_0, A0, A1);
NANDC2x1 inst_and_b3_1_0 ( imd_Y3, wire3_0_0, wire3_0_1);
NANDC2x1 inst_and_b2_0_0 ( imd_wire2_0_0, A0_inv, A1);
NANDC2x1 inst_clockedAND_b2_2 ( imd_YF2, CLK, Y2);
NANDC2x1 inst_and_b2_0_1 ( imd_wire2_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b2_1_0 ( imd_Y2, wire2_0_0, wire2_0_1);
NANDC2x1 inst_and_b1_0_0 ( imd_wire1_0_0, A0, A1_inv);
NANDC2x1 inst_clockedAND_b1_1 ( imd_YF1, CLK, Y1);
NANDC2x1 inst_and_b1_0_1 ( imd_wire1_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b1_1_0 ( imd_Y1, wire1_0_0, wire1_0_1);
NANDC2x1 inst_and_b0_0_0 ( imd_wire0_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b0_0_1 ( imd_wire0_0_1, A2_inv, A3_inv);
NANDC2x1 inst_clockedAND_b0_0 ( imd_YF0, CLK, Y0);
NANDC2x1 inst_and_b0_1_0 ( imd_Y0, wire0_0_0, wire0_0_1);
INVC inst_clockedinv_b15_15 ( YF15, imd_YF15);
INVC inst_inv_b15_1_0 ( Y15, imd_Y15);
INVC inst_inv_b15_0_1 ( wire15_0_1, imd_wire15_0_1);
INVC inst_inv_b15_0_0 ( wire15_0_0, imd_wire15_0_0);
INVC inst_clockedinv_b14_14 ( YF14, imd_YF14);
INVC inst_inv_b14_1_0 ( Y14, imd_Y14);
INVC inst_inv_b14_0_1 ( wire14_0_1, imd_wire14_0_1);
INVC inst_inv_b14_0_0 ( wire14_0_0, imd_wire14_0_0);
INVC inst_clockedinv_b13_13 ( YF13, imd_YF13);
INVC inst_inv_b13_1_0 ( Y13, imd_Y13);
INVC inst_inv_b13_0_1 ( wire13_0_1, imd_wire13_0_1);
INVC inst_inv_b13_0_0 ( wire13_0_0, imd_wire13_0_0);
INVC inst_clockedinv_b12_12 ( YF12, imd_YF12);
INVC inst_inv_b12_1_0 ( Y12, imd_Y12);
INVC inst_inv_b12_0_1 ( wire12_0_1, imd_wire12_0_1);
INVC inst_inv_b12_0_0 ( wire12_0_0, imd_wire12_0_0);
INVC inst_clockedinv_b11_11 ( YF11, imd_YF11);
INVC inst_inv_b11_1_0 ( Y11, imd_Y11);
INVC inst_inv_b11_0_1 ( wire11_0_1, imd_wire11_0_1);
INVC inst_inv_b11_0_0 ( wire11_0_0, imd_wire11_0_0);
INVC inst_clockedinv_b10_10 ( YF10, imd_YF10);
INVC inst_inv_b10_1_0 ( Y10, imd_Y10);
INVC inst_inv_b10_0_1 ( wire10_0_1, imd_wire10_0_1);
INVC inst_inv_b10_0_0 ( wire10_0_0, imd_wire10_0_0);
INVC inst_clockedinv_b9_9 ( YF9, imd_YF9);
INVC inst_inv_b9_1_0 ( Y9, imd_Y9);
INVC inst_inv_b9_0_1 ( wire9_0_1, imd_wire9_0_1);
INVC inst_inv_b9_0_0 ( wire9_0_0, imd_wire9_0_0);
INVC inst_inv_b8_0_1 ( wire8_0_1, imd_wire8_0_1);
INVC inst_inv_b8_1_0 ( Y8, imd_Y8);
INVC inst_clockedinv_b8_8 ( YF8, imd_YF8);
INVC inst_inv_b8_0_0 ( wire8_0_0, imd_wire8_0_0);
INVC inst_clockedinv_b7_7 ( YF7, imd_YF7);
INVC inst_inv_b7_1_0 ( Y7, imd_Y7);
INVC inst_inv_b7_0_1 ( wire7_0_1, imd_wire7_0_1);
INVC inst_inv_b7_0_0 ( wire7_0_0, imd_wire7_0_0);
INVC inst_clockedinv_b6_6 ( YF6, imd_YF6);
INVC inst_inv_b6_1_0 ( Y6, imd_Y6);
INVC inst_inv_b6_0_1 ( wire6_0_1, imd_wire6_0_1);
INVC inst_inv_b6_0_0 ( wire6_0_0, imd_wire6_0_0);
INVC inst_clockedinv_b5_5 ( YF5, imd_YF5);
INVC inst_inv_b5_1_0 ( Y5, imd_Y5);
INVC inst_inv_b5_0_1 ( wire5_0_1, imd_wire5_0_1);
INVC inst_inv_b5_0_0 ( wire5_0_0, imd_wire5_0_0);
INVC inst_inv_b4_0_1 ( wire4_0_1, imd_wire4_0_1);
INVC inst_inv_b4_1_0 ( Y4, imd_Y4);
INVC inst_clockedinv_b4_4 ( YF4, imd_YF4);
INVC inst_inv_b4_0_0 ( wire4_0_0, imd_wire4_0_0);
INVC inst_clockedinv_b3_3 ( YF3, imd_YF3);
INVC inst_inv_b3_1_0 ( Y3, imd_Y3);
INVC inst_inv_b3_0_1 ( wire3_0_1, imd_wire3_0_1);
INVC inst_inv_b3_0_0 ( wire3_0_0, imd_wire3_0_0);
INVC inst_inv_b2_0_0 ( wire2_0_0, imd_wire2_0_0);
INVC inst_inv_b2_1_0 ( Y2, imd_Y2);
INVC inst_clockedinv_b2_2 ( YF2, imd_YF2);
INVC inst_inv_b2_0_1 ( wire2_0_1, imd_wire2_0_1);
INVC inst_inv_b1_0_0 ( wire1_0_0, imd_wire1_0_0);
INVC inst_inv_b1_1_0 ( Y1, imd_Y1);
INVC inst_clockedinv_b1_1 ( YF1, imd_YF1);
INVC inst_inv_b1_0_1 ( wire1_0_1, imd_wire1_0_1);
INVC inst_inv_b0_0_0 ( wire0_0_0, imd_wire0_0_0);
INVC inst_inv_b0_0_1 ( wire0_0_1, imd_wire0_0_1);
INVC inst_inv_b0_1_0 ( Y0, imd_Y0);
INVC inst_clockedinv_b0_0 ( YF0, imd_YF0);

endmodule
// Library - sram_compiled_r128_c128_w8, Cell - invCol, View -
//schematic
// LAST TIME SAVED: Apr 20 20:07:34 2021
// NETLIST TIME: Apr 21 18:57:09 2021
`timescale 1ns / 1ps 

module invCol ( A0, A1, A2, A3, Abar0, Abar1, Abar2, Abar3 );

output  Abar0, Abar1, Abar2, Abar3;

input  A0, A1, A2, A3;


specify 
    specparam CDS_LIBNAME  = "sram_compiled_r128_c128_w8";
    specparam CDS_CELLNAME = "invCol";
    specparam CDS_VIEWNAME = "schematic";
endspecify

INVD wire3 ( Abar3, A3);
INVD wire2 ( Abar2, A2);
INVD wire1 ( Abar1, A1);
INVD wire0 ( Abar0, A0);

endmodule
// Library - sram_compiled_r128_c128_w8, Cell - columnMux, View -
//schematic
// LAST TIME SAVED: Apr 20 20:07:34 2021
// NETLIST TIME: Apr 21 18:57:09 2021
`timescale 1ns / 1ps 

module columnMux ( A0, Abar0, A1, Abar1, A2, Abar2, A3, Abar3, A4,
     Abar4, A5, Abar5, A6, Abar6, A7, Abar7, A8, Abar8, A9, Abar9, A10,
     Abar10, A11, Abar11, A12, Abar12, A13, Abar13, A14, Abar14, A15,
     Abar15, sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8,
     sel9, sel10, sel11, sel12, sel13, sel14, sel15, Y, Ybar );

output  Y, Ybar;

input  A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14,
     A15, Abar0, Abar1, Abar2, Abar3, Abar4, Abar5, Abar6, Abar7,
     Abar8, Abar9, Abar10, Abar11, Abar12, Abar13, Abar14, Abar15,
     sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8, sel9, sel10,
     sel11, sel12, sel13, sel14, sel15;


specify 
    specparam CDS_LIBNAME  = "sram_compiled_r128_c128_w8";
    specparam CDS_CELLNAME = "columnMux";
    specparam CDS_VIEWNAME = "schematic";
endspecify

muxTrans wire31 ( Abar15, Ybar, sel15);
muxTrans wire30 ( A15, Y, sel15);
muxTrans wire29 ( Abar14, Ybar, sel14);
muxTrans wire28 ( A14, Y, sel14);
muxTrans wire27 ( Abar13, Ybar, sel13);
muxTrans wire26 ( A13, Y, sel13);
muxTrans wire25 ( Abar12, Ybar, sel12);
muxTrans wire24 ( A12, Y, sel12);
muxTrans wire23 ( Abar11, Ybar, sel11);
muxTrans wire22 ( A11, Y, sel11);
muxTrans wire21 ( Abar10, Ybar, sel10);
muxTrans wire20 ( A10, Y, sel10);
muxTrans wire19 ( Abar9, Ybar, sel9);
muxTrans wire18 ( A9, Y, sel9);
muxTrans wire17 ( Abar8, Ybar, sel8);
muxTrans wire16 ( A8, Y, sel8);
muxTrans wire15 ( Abar7, Ybar, sel7);
muxTrans wire14 ( A7, Y, sel7);
muxTrans wire13 ( Abar6, Ybar, sel6);
muxTrans wire12 ( A6, Y, sel6);
muxTrans wire11 ( Abar5, Ybar, sel5);
muxTrans wire10 ( A5, Y, sel5);
muxTrans wire9 ( Abar4, Ybar, sel4);
muxTrans wire8 ( A4, Y, sel4);
muxTrans wire7 ( Abar3, Ybar, sel3);
muxTrans wire6 ( A3, Y, sel3);
muxTrans wire5 ( Abar2, Ybar, sel2);
muxTrans wire4 ( A2, Y, sel2);
muxTrans wire3 ( Abar1, Ybar, sel1);
muxTrans wire2 ( A1, Y, sel1);
muxTrans wire1 ( Abar0, Ybar, sel0);
muxTrans wire0 ( A0, Y, sel0);

endmodule
// Library - sram_compiled_r128_c128_w8, Cell - invRow, View -
//schematic
// LAST TIME SAVED: Apr 20 20:07:34 2021
// NETLIST TIME: Apr 21 18:57:09 2021
`timescale 1ns / 1ps 

module invRow ( A0, A1, A2, A3, A4, A5, A6, Abar0, Abar1, Abar2, Abar3,
     Abar4, Abar5, Abar6 );

output  Abar0, Abar1, Abar2, Abar3, Abar4, Abar5, Abar6;

input  A0, A1, A2, A3, A4, A5, A6;


specify 
    specparam CDS_LIBNAME  = "sram_compiled_r128_c128_w8";
    specparam CDS_CELLNAME = "invRow";
    specparam CDS_VIEWNAME = "schematic";
endspecify

INVD wire6 ( Abar6, A6);
INVD wire5 ( Abar5, A5);
INVD wire4 ( Abar4, A4);
INVD wire3 ( Abar3, A3);
INVD wire2 ( Abar2, A2);
INVD wire1 ( Abar1, A1);
INVD wire0 ( Abar0, A0);

endmodule
// Library - sram_compiled_r128_c128_w8, Cell - rowDecoder, View -
//schematic
// LAST TIME SAVED: Apr 20 20:07:34 2021
// NETLIST TIME: Apr 21 18:57:10 2021
`timescale 1ns / 1ps 

module rowDecoder ( A0, A0_inv, A1, A1_inv, A2, A2_inv, A3, A3_inv, A4,
     A4_inv, A5, A5_inv, A6, A6_inv, CLK, YF0, YF1, YF2, YF3, YF4, YF5,
     YF6, YF7, YF8, YF9, YF10, YF11, YF12, YF13, YF14, YF15, YF16,
     YF17, YF18, YF19, YF20, YF21, YF22, YF23, YF24, YF25, YF26, YF27,
     YF28, YF29, YF30, YF31, YF32, YF33, YF34, YF35, YF36, YF37, YF38,
     YF39, YF40, YF41, YF42, YF43, YF44, YF45, YF46, YF47, YF48, YF49,
     YF50, YF51, YF52, YF53, YF54, YF55, YF56, YF57, YF58, YF59, YF60,
     YF61, YF62, YF63, YF64, YF65, YF66, YF67, YF68, YF69, YF70, YF71,
     YF72, YF73, YF74, YF75, YF76, YF77, YF78, YF79, YF80, YF81, YF82,
     YF83, YF84, YF85, YF86, YF87, YF88, YF89, YF90, YF91, YF92, YF93,
     YF94, YF95, YF96, YF97, YF98, YF99, YF100, YF101, YF102, YF103,
     YF104, YF105, YF106, YF107, YF108, YF109, YF110, YF111, YF112,
     YF113, YF114, YF115, YF116, YF117, YF118, YF119, YF120, YF121,
     YF122, YF123, YF124, YF125, YF126, YF127 );

output  YF0, YF1, YF2, YF3, YF4, YF5, YF6, YF7, YF8, YF9, YF10, YF11,
     YF12, YF13, YF14, YF15, YF16, YF17, YF18, YF19, YF20, YF21, YF22,
     YF23, YF24, YF25, YF26, YF27, YF28, YF29, YF30, YF31, YF32, YF33,
     YF34, YF35, YF36, YF37, YF38, YF39, YF40, YF41, YF42, YF43, YF44,
     YF45, YF46, YF47, YF48, YF49, YF50, YF51, YF52, YF53, YF54, YF55,
     YF56, YF57, YF58, YF59, YF60, YF61, YF62, YF63, YF64, YF65, YF66,
     YF67, YF68, YF69, YF70, YF71, YF72, YF73, YF74, YF75, YF76, YF77,
     YF78, YF79, YF80, YF81, YF82, YF83, YF84, YF85, YF86, YF87, YF88,
     YF89, YF90, YF91, YF92, YF93, YF94, YF95, YF96, YF97, YF98, YF99,
     YF100, YF101, YF102, YF103, YF104, YF105, YF106, YF107, YF108,
     YF109, YF110, YF111, YF112, YF113, YF114, YF115, YF116, YF117,
     YF118, YF119, YF120, YF121, YF122, YF123, YF124, YF125, YF126,
     YF127;

input  A0, A0_inv, A1, A1_inv, A2, A2_inv, A3, A3_inv, A4, A4_inv, A5,
     A5_inv, A6, A6_inv, CLK;


specify 
    specparam CDS_LIBNAME  = "sram_compiled_r128_c128_w8";
    specparam CDS_CELLNAME = "rowDecoder";
    specparam CDS_VIEWNAME = "schematic";
endspecify

NANDC2x1 inst_clockedAND_b127_127 ( imd_YF127, CLK, Y127);
NANDC2x1 inst_and_b127_1_1 ( imd_wire127_1_1, A6, wire127_0_2);
NANDC2x1 inst_and_b127_0_2 ( imd_wire127_0_2, A4, A5);
NANDC2x1 inst_and_b127_2_0 ( imd_Y127, wire127_1_0, wire127_1_1);
NANDC2x1 inst_and_b127_0_1 ( imd_wire127_0_1, A2, A3);
NANDC2x1 inst_and_b127_0_0 ( imd_wire127_0_0, A0, A1);
NANDC2x1 inst_and_b127_1_0 ( imd_wire127_1_0, wire127_0_0,
     wire127_0_1);
NANDC2x1 inst_clockedAND_b126_126 ( imd_YF126, CLK, Y126);
NANDC2x1 inst_and_b126_1_1 ( imd_wire126_1_1, A6, wire126_0_2);
NANDC2x1 inst_and_b126_0_2 ( imd_wire126_0_2, A4, A5);
NANDC2x1 inst_and_b126_2_0 ( imd_Y126, wire126_1_0, wire126_1_1);
NANDC2x1 inst_and_b126_0_1 ( imd_wire126_0_1, A2, A3);
NANDC2x1 inst_and_b126_0_0 ( imd_wire126_0_0, A0_inv, A1);
NANDC2x1 inst_and_b126_1_0 ( imd_wire126_1_0, wire126_0_0,
     wire126_0_1);
NANDC2x1 inst_clockedAND_b125_125 ( imd_YF125, CLK, Y125);
NANDC2x1 inst_and_b125_1_1 ( imd_wire125_1_1, A6, wire125_0_2);
NANDC2x1 inst_and_b125_0_2 ( imd_wire125_0_2, A4, A5);
NANDC2x1 inst_and_b125_2_0 ( imd_Y125, wire125_1_0, wire125_1_1);
NANDC2x1 inst_and_b125_0_1 ( imd_wire125_0_1, A2, A3);
NANDC2x1 inst_and_b125_0_0 ( imd_wire125_0_0, A0, A1_inv);
NANDC2x1 inst_and_b125_1_0 ( imd_wire125_1_0, wire125_0_0,
     wire125_0_1);
NANDC2x1 inst_clockedAND_b124_124 ( imd_YF124, CLK, Y124);
NANDC2x1 inst_and_b124_1_1 ( imd_wire124_1_1, A6, wire124_0_2);
NANDC2x1 inst_and_b124_0_2 ( imd_wire124_0_2, A4, A5);
NANDC2x1 inst_and_b124_2_0 ( imd_Y124, wire124_1_0, wire124_1_1);
NANDC2x1 inst_and_b124_0_1 ( imd_wire124_0_1, A2, A3);
NANDC2x1 inst_and_b124_0_0 ( imd_wire124_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b124_1_0 ( imd_wire124_1_0, wire124_0_0,
     wire124_0_1);
NANDC2x1 inst_clockedAND_b123_123 ( imd_YF123, CLK, Y123);
NANDC2x1 inst_and_b123_1_1 ( imd_wire123_1_1, A6, wire123_0_2);
NANDC2x1 inst_and_b123_0_2 ( imd_wire123_0_2, A4, A5);
NANDC2x1 inst_and_b123_2_0 ( imd_Y123, wire123_1_0, wire123_1_1);
NANDC2x1 inst_and_b123_0_1 ( imd_wire123_0_1, A2_inv, A3);
NANDC2x1 inst_and_b123_0_0 ( imd_wire123_0_0, A0, A1);
NANDC2x1 inst_and_b123_1_0 ( imd_wire123_1_0, wire123_0_0,
     wire123_0_1);
NANDC2x1 inst_clockedAND_b122_122 ( imd_YF122, CLK, Y122);
NANDC2x1 inst_and_b122_1_1 ( imd_wire122_1_1, A6, wire122_0_2);
NANDC2x1 inst_and_b122_0_2 ( imd_wire122_0_2, A4, A5);
NANDC2x1 inst_and_b122_2_0 ( imd_Y122, wire122_1_0, wire122_1_1);
NANDC2x1 inst_and_b122_0_1 ( imd_wire122_0_1, A2_inv, A3);
NANDC2x1 inst_and_b122_0_0 ( imd_wire122_0_0, A0_inv, A1);
NANDC2x1 inst_and_b122_1_0 ( imd_wire122_1_0, wire122_0_0,
     wire122_0_1);
NANDC2x1 inst_clockedAND_b121_121 ( imd_YF121, CLK, Y121);
NANDC2x1 inst_and_b121_1_1 ( imd_wire121_1_1, A6, wire121_0_2);
NANDC2x1 inst_and_b121_0_2 ( imd_wire121_0_2, A4, A5);
NANDC2x1 inst_and_b121_2_0 ( imd_Y121, wire121_1_0, wire121_1_1);
NANDC2x1 inst_and_b121_0_1 ( imd_wire121_0_1, A2_inv, A3);
NANDC2x1 inst_and_b121_0_0 ( imd_wire121_0_0, A0, A1_inv);
NANDC2x1 inst_and_b121_1_0 ( imd_wire121_1_0, wire121_0_0,
     wire121_0_1);
NANDC2x1 inst_clockedAND_b120_120 ( imd_YF120, CLK, Y120);
NANDC2x1 inst_and_b120_1_1 ( imd_wire120_1_1, A6, wire120_0_2);
NANDC2x1 inst_and_b120_0_2 ( imd_wire120_0_2, A4, A5);
NANDC2x1 inst_and_b120_2_0 ( imd_Y120, wire120_1_0, wire120_1_1);
NANDC2x1 inst_and_b120_0_1 ( imd_wire120_0_1, A2_inv, A3);
NANDC2x1 inst_and_b120_0_0 ( imd_wire120_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b120_1_0 ( imd_wire120_1_0, wire120_0_0,
     wire120_0_1);
NANDC2x1 inst_clockedAND_b119_119 ( imd_YF119, CLK, Y119);
NANDC2x1 inst_and_b119_1_1 ( imd_wire119_1_1, A6, wire119_0_2);
NANDC2x1 inst_and_b119_0_2 ( imd_wire119_0_2, A4, A5);
NANDC2x1 inst_and_b119_2_0 ( imd_Y119, wire119_1_0, wire119_1_1);
NANDC2x1 inst_and_b119_0_1 ( imd_wire119_0_1, A2, A3_inv);
NANDC2x1 inst_and_b119_0_0 ( imd_wire119_0_0, A0, A1);
NANDC2x1 inst_and_b119_1_0 ( imd_wire119_1_0, wire119_0_0,
     wire119_0_1);
NANDC2x1 inst_clockedAND_b118_118 ( imd_YF118, CLK, Y118);
NANDC2x1 inst_and_b118_1_1 ( imd_wire118_1_1, A6, wire118_0_2);
NANDC2x1 inst_and_b118_0_2 ( imd_wire118_0_2, A4, A5);
NANDC2x1 inst_and_b118_2_0 ( imd_Y118, wire118_1_0, wire118_1_1);
NANDC2x1 inst_and_b118_0_1 ( imd_wire118_0_1, A2, A3_inv);
NANDC2x1 inst_and_b118_0_0 ( imd_wire118_0_0, A0_inv, A1);
NANDC2x1 inst_and_b118_1_0 ( imd_wire118_1_0, wire118_0_0,
     wire118_0_1);
NANDC2x1 inst_clockedAND_b117_117 ( imd_YF117, CLK, Y117);
NANDC2x1 inst_and_b117_1_1 ( imd_wire117_1_1, A6, wire117_0_2);
NANDC2x1 inst_and_b117_0_2 ( imd_wire117_0_2, A4, A5);
NANDC2x1 inst_and_b117_2_0 ( imd_Y117, wire117_1_0, wire117_1_1);
NANDC2x1 inst_and_b117_0_1 ( imd_wire117_0_1, A2, A3_inv);
NANDC2x1 inst_and_b117_0_0 ( imd_wire117_0_0, A0, A1_inv);
NANDC2x1 inst_and_b117_1_0 ( imd_wire117_1_0, wire117_0_0,
     wire117_0_1);
NANDC2x1 inst_clockedAND_b116_116 ( imd_YF116, CLK, Y116);
NANDC2x1 inst_and_b116_1_1 ( imd_wire116_1_1, A6, wire116_0_2);
NANDC2x1 inst_and_b116_0_2 ( imd_wire116_0_2, A4, A5);
NANDC2x1 inst_and_b116_2_0 ( imd_Y116, wire116_1_0, wire116_1_1);
NANDC2x1 inst_and_b116_0_1 ( imd_wire116_0_1, A2, A3_inv);
NANDC2x1 inst_and_b116_0_0 ( imd_wire116_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b116_1_0 ( imd_wire116_1_0, wire116_0_0,
     wire116_0_1);
NANDC2x1 inst_clockedAND_b115_115 ( imd_YF115, CLK, Y115);
NANDC2x1 inst_and_b115_1_1 ( imd_wire115_1_1, A6, wire115_0_2);
NANDC2x1 inst_and_b115_0_2 ( imd_wire115_0_2, A4, A5);
NANDC2x1 inst_and_b115_2_0 ( imd_Y115, wire115_1_0, wire115_1_1);
NANDC2x1 inst_and_b115_0_1 ( imd_wire115_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b115_0_0 ( imd_wire115_0_0, A0, A1);
NANDC2x1 inst_and_b115_1_0 ( imd_wire115_1_0, wire115_0_0,
     wire115_0_1);
NANDC2x1 inst_clockedAND_b114_114 ( imd_YF114, CLK, Y114);
NANDC2x1 inst_and_b114_1_1 ( imd_wire114_1_1, A6, wire114_0_2);
NANDC2x1 inst_and_b114_0_2 ( imd_wire114_0_2, A4, A5);
NANDC2x1 inst_and_b114_2_0 ( imd_Y114, wire114_1_0, wire114_1_1);
NANDC2x1 inst_and_b114_0_1 ( imd_wire114_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b114_0_0 ( imd_wire114_0_0, A0_inv, A1);
NANDC2x1 inst_and_b114_1_0 ( imd_wire114_1_0, wire114_0_0,
     wire114_0_1);
NANDC2x1 inst_clockedAND_b113_113 ( imd_YF113, CLK, Y113);
NANDC2x1 inst_and_b113_1_1 ( imd_wire113_1_1, A6, wire113_0_2);
NANDC2x1 inst_and_b113_0_2 ( imd_wire113_0_2, A4, A5);
NANDC2x1 inst_and_b113_2_0 ( imd_Y113, wire113_1_0, wire113_1_1);
NANDC2x1 inst_and_b113_0_1 ( imd_wire113_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b113_0_0 ( imd_wire113_0_0, A0, A1_inv);
NANDC2x1 inst_and_b113_1_0 ( imd_wire113_1_0, wire113_0_0,
     wire113_0_1);
NANDC2x1 inst_clockedAND_b112_112 ( imd_YF112, CLK, Y112);
NANDC2x1 inst_and_b112_1_1 ( imd_wire112_1_1, A6, wire112_0_2);
NANDC2x1 inst_and_b112_0_2 ( imd_wire112_0_2, A4, A5);
NANDC2x1 inst_and_b112_2_0 ( imd_Y112, wire112_1_0, wire112_1_1);
NANDC2x1 inst_and_b112_0_1 ( imd_wire112_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b112_0_0 ( imd_wire112_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b112_1_0 ( imd_wire112_1_0, wire112_0_0,
     wire112_0_1);
NANDC2x1 inst_and_b111_0_1 ( imd_wire111_0_1, A2, A3);
NANDC2x1 inst_and_b110_0_1 ( imd_wire110_0_1, A2, A3);
NANDC2x1 inst_and_b111_0_0 ( imd_wire111_0_0, A0, A1);
NANDC2x1 inst_and_b111_1_0 ( imd_wire111_1_0, wire111_0_0,
     wire111_0_1);
NANDC2x1 inst_clockedAND_b110_110 ( imd_YF110, CLK, Y110);
NANDC2x1 inst_and_b110_1_1 ( imd_wire110_1_1, A6, wire110_0_2);
NANDC2x1 inst_and_b110_1_0 ( imd_wire110_1_0, wire110_0_0,
     wire110_0_1);
NANDC2x1 inst_and_b110_0_0 ( imd_wire110_0_0, A0_inv, A1);
NANDC2x1 inst_and_b110_2_0 ( imd_Y110, wire110_1_0, wire110_1_1);
NANDC2x1 inst_clockedAND_b111_111 ( imd_YF111, CLK, Y111);
NANDC2x1 inst_and_b111_2_0 ( imd_Y111, wire111_1_0, wire111_1_1);
NANDC2x1 inst_and_b111_1_1 ( imd_wire111_1_1, A6, wire111_0_2);
NANDC2x1 inst_and_b111_0_2 ( imd_wire111_0_2, A4_inv, A5);
NANDC2x1 inst_and_b110_0_2 ( imd_wire110_0_2, A4_inv, A5);
NANDC2x1 inst_clockedAND_b109_109 ( imd_YF109, CLK, Y109);
NANDC2x1 inst_and_b109_1_1 ( imd_wire109_1_1, A6, wire109_0_2);
NANDC2x1 inst_and_b109_0_2 ( imd_wire109_0_2, A4_inv, A5);
NANDC2x1 inst_and_b109_2_0 ( imd_Y109, wire109_1_0, wire109_1_1);
NANDC2x1 inst_and_b109_0_1 ( imd_wire109_0_1, A2, A3);
NANDC2x1 inst_and_b109_0_0 ( imd_wire109_0_0, A0, A1_inv);
NANDC2x1 inst_and_b109_1_0 ( imd_wire109_1_0, wire109_0_0,
     wire109_0_1);
NANDC2x1 inst_clockedAND_b108_108 ( imd_YF108, CLK, Y108);
NANDC2x1 inst_and_b108_1_1 ( imd_wire108_1_1, A6, wire108_0_2);
NANDC2x1 inst_and_b108_0_2 ( imd_wire108_0_2, A4_inv, A5);
NANDC2x1 inst_and_b108_2_0 ( imd_Y108, wire108_1_0, wire108_1_1);
NANDC2x1 inst_and_b108_0_1 ( imd_wire108_0_1, A2, A3);
NANDC2x1 inst_and_b108_0_0 ( imd_wire108_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b108_1_0 ( imd_wire108_1_0, wire108_0_0,
     wire108_0_1);
NANDC2x1 inst_clockedAND_b107_107 ( imd_YF107, CLK, Y107);
NANDC2x1 inst_and_b107_1_1 ( imd_wire107_1_1, A6, wire107_0_2);
NANDC2x1 inst_and_b107_0_2 ( imd_wire107_0_2, A4_inv, A5);
NANDC2x1 inst_and_b107_2_0 ( imd_Y107, wire107_1_0, wire107_1_1);
NANDC2x1 inst_and_b107_0_1 ( imd_wire107_0_1, A2_inv, A3);
NANDC2x1 inst_and_b107_0_0 ( imd_wire107_0_0, A0, A1);
NANDC2x1 inst_and_b107_1_0 ( imd_wire107_1_0, wire107_0_0,
     wire107_0_1);
NANDC2x1 inst_clockedAND_b106_106 ( imd_YF106, CLK, Y106);
NANDC2x1 inst_and_b106_1_1 ( imd_wire106_1_1, A6, wire106_0_2);
NANDC2x1 inst_and_b106_0_2 ( imd_wire106_0_2, A4_inv, A5);
NANDC2x1 inst_and_b106_2_0 ( imd_Y106, wire106_1_0, wire106_1_1);
NANDC2x1 inst_and_b106_0_1 ( imd_wire106_0_1, A2_inv, A3);
NANDC2x1 inst_and_b106_0_0 ( imd_wire106_0_0, A0_inv, A1);
NANDC2x1 inst_and_b106_1_0 ( imd_wire106_1_0, wire106_0_0,
     wire106_0_1);
NANDC2x1 inst_clockedAND_b105_105 ( imd_YF105, CLK, Y105);
NANDC2x1 inst_and_b105_1_1 ( imd_wire105_1_1, A6, wire105_0_2);
NANDC2x1 inst_and_b105_0_2 ( imd_wire105_0_2, A4_inv, A5);
NANDC2x1 inst_and_b105_2_0 ( imd_Y105, wire105_1_0, wire105_1_1);
NANDC2x1 inst_and_b105_0_1 ( imd_wire105_0_1, A2_inv, A3);
NANDC2x1 inst_and_b105_0_0 ( imd_wire105_0_0, A0, A1_inv);
NANDC2x1 inst_and_b105_1_0 ( imd_wire105_1_0, wire105_0_0,
     wire105_0_1);
NANDC2x1 inst_clockedAND_b104_104 ( imd_YF104, CLK, Y104);
NANDC2x1 inst_and_b104_1_1 ( imd_wire104_1_1, A6, wire104_0_2);
NANDC2x1 inst_and_b104_0_2 ( imd_wire104_0_2, A4_inv, A5);
NANDC2x1 inst_and_b104_2_0 ( imd_Y104, wire104_1_0, wire104_1_1);
NANDC2x1 inst_and_b104_0_1 ( imd_wire104_0_1, A2_inv, A3);
NANDC2x1 inst_and_b104_0_0 ( imd_wire104_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b104_1_0 ( imd_wire104_1_0, wire104_0_0,
     wire104_0_1);
NANDC2x1 inst_clockedAND_b103_103 ( imd_YF103, CLK, Y103);
NANDC2x1 inst_and_b103_1_1 ( imd_wire103_1_1, A6, wire103_0_2);
NANDC2x1 inst_and_b103_0_2 ( imd_wire103_0_2, A4_inv, A5);
NANDC2x1 inst_and_b103_2_0 ( imd_Y103, wire103_1_0, wire103_1_1);
NANDC2x1 inst_and_b103_0_1 ( imd_wire103_0_1, A2, A3_inv);
NANDC2x1 inst_and_b103_0_0 ( imd_wire103_0_0, A0, A1);
NANDC2x1 inst_and_b103_1_0 ( imd_wire103_1_0, wire103_0_0,
     wire103_0_1);
NANDC2x1 inst_clockedAND_b102_102 ( imd_YF102, CLK, Y102);
NANDC2x1 inst_and_b102_1_1 ( imd_wire102_1_1, A6, wire102_0_2);
NANDC2x1 inst_and_b102_0_2 ( imd_wire102_0_2, A4_inv, A5);
NANDC2x1 inst_and_b102_2_0 ( imd_Y102, wire102_1_0, wire102_1_1);
NANDC2x1 inst_and_b102_0_1 ( imd_wire102_0_1, A2, A3_inv);
NANDC2x1 inst_and_b102_0_0 ( imd_wire102_0_0, A0_inv, A1);
NANDC2x1 inst_and_b102_1_0 ( imd_wire102_1_0, wire102_0_0,
     wire102_0_1);
NANDC2x1 inst_clockedAND_b101_101 ( imd_YF101, CLK, Y101);
NANDC2x1 inst_and_b101_1_1 ( imd_wire101_1_1, A6, wire101_0_2);
NANDC2x1 inst_and_b101_0_2 ( imd_wire101_0_2, A4_inv, A5);
NANDC2x1 inst_and_b101_2_0 ( imd_Y101, wire101_1_0, wire101_1_1);
NANDC2x1 inst_and_b101_0_1 ( imd_wire101_0_1, A2, A3_inv);
NANDC2x1 inst_and_b101_0_0 ( imd_wire101_0_0, A0, A1_inv);
NANDC2x1 inst_and_b101_1_0 ( imd_wire101_1_0, wire101_0_0,
     wire101_0_1);
NANDC2x1 inst_clockedAND_b100_100 ( imd_YF100, CLK, Y100);
NANDC2x1 inst_and_b100_2_0 ( imd_Y100, wire100_1_0, wire100_1_1);
NANDC2x1 inst_and_b100_0_1 ( imd_wire100_0_1, A2, A3_inv);
NANDC2x1 inst_and_b100_0_0 ( imd_wire100_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b100_1_0 ( imd_wire100_1_0, wire100_0_0,
     wire100_0_1);
NANDC2x1 inst_clockedAND_b99_99 ( imd_YF99, CLK, Y99);
NANDC2x1 inst_and_b99_1_1 ( imd_wire99_1_1, A6, wire99_0_2);
NANDC2x1 inst_and_b99_0_2 ( imd_wire99_0_2, A4_inv, A5);
NANDC2x1 inst_and_b99_2_0 ( imd_Y99, wire99_1_0, wire99_1_1);
NANDC2x1 inst_and_b99_0_1 ( imd_wire99_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b99_0_0 ( imd_wire99_0_0, A0, A1);
NANDC2x1 inst_and_b99_1_0 ( imd_wire99_1_0, wire99_0_0, wire99_0_1);
NANDC2x1 inst_clockedAND_b98_98 ( imd_YF98, CLK, Y98);
NANDC2x1 inst_and_b98_1_1 ( imd_wire98_1_1, A6, wire98_0_2);
NANDC2x1 inst_and_b98_0_2 ( imd_wire98_0_2, A4_inv, A5);
NANDC2x1 inst_and_b98_2_0 ( imd_Y98, wire98_1_0, wire98_1_1);
NANDC2x1 inst_and_b98_0_1 ( imd_wire98_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b98_0_0 ( imd_wire98_0_0, A0_inv, A1);
NANDC2x1 inst_and_b98_1_0 ( imd_wire98_1_0, wire98_0_0, wire98_0_1);
NANDC2x1 inst_clockedAND_b97_97 ( imd_YF97, CLK, Y97);
NANDC2x1 inst_and_b97_1_1 ( imd_wire97_1_1, A6, wire97_0_2);
NANDC2x1 inst_and_b97_0_2 ( imd_wire97_0_2, A4_inv, A5);
NANDC2x1 inst_and_b97_2_0 ( imd_Y97, wire97_1_0, wire97_1_1);
NANDC2x1 inst_and_b97_0_1 ( imd_wire97_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b97_0_0 ( imd_wire97_0_0, A0, A1_inv);
NANDC2x1 inst_and_b97_1_0 ( imd_wire97_1_0, wire97_0_0, wire97_0_1);
NANDC2x1 inst_clockedAND_b96_96 ( imd_YF96, CLK, Y96);
NANDC2x1 inst_and_b96_1_1 ( imd_wire96_1_1, A6, wire96_0_2);
NANDC2x1 inst_and_b96_0_2 ( imd_wire96_0_2, A4_inv, A5);
NANDC2x1 inst_and_b96_2_0 ( imd_Y96, wire96_1_0, wire96_1_1);
NANDC2x1 inst_and_b96_0_1 ( imd_wire96_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b96_0_0 ( imd_wire96_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b96_1_0 ( imd_wire96_1_0, wire96_0_0, wire96_0_1);
NANDC2x1 inst_clockedAND_b95_95 ( imd_YF95, CLK, Y95);
NANDC2x1 inst_and_b95_1_1 ( imd_wire95_1_1, A6, wire95_0_2);
NANDC2x1 inst_and_b95_0_2 ( imd_wire95_0_2, A4, A5_inv);
NANDC2x1 inst_and_b95_2_0 ( imd_Y95, wire95_1_0, wire95_1_1);
NANDC2x1 inst_and_b95_0_1 ( imd_wire95_0_1, A2, A3);
NANDC2x1 inst_and_b95_0_0 ( imd_wire95_0_0, A0, A1);
NANDC2x1 inst_and_b95_1_0 ( imd_wire95_1_0, wire95_0_0, wire95_0_1);
NANDC2x1 inst_clockedAND_b94_94 ( imd_YF94, CLK, Y94);
NANDC2x1 inst_and_b94_1_1 ( imd_wire94_1_1, A6, wire94_0_2);
NANDC2x1 inst_and_b94_0_2 ( imd_wire94_0_2, A4, A5_inv);
NANDC2x1 inst_and_b94_2_0 ( imd_Y94, wire94_1_0, wire94_1_1);
NANDC2x1 inst_and_b94_0_1 ( imd_wire94_0_1, A2, A3);
NANDC2x1 inst_and_b94_0_0 ( imd_wire94_0_0, A0_inv, A1);
NANDC2x1 inst_and_b94_1_0 ( imd_wire94_1_0, wire94_0_0, wire94_0_1);
NANDC2x1 inst_clockedAND_b93_93 ( imd_YF93, CLK, Y93);
NANDC2x1 inst_and_b93_1_1 ( imd_wire93_1_1, A6, wire93_0_2);
NANDC2x1 inst_and_b93_0_2 ( imd_wire93_0_2, A4, A5_inv);
NANDC2x1 inst_and_b93_2_0 ( imd_Y93, wire93_1_0, wire93_1_1);
NANDC2x1 inst_and_b93_0_1 ( imd_wire93_0_1, A2, A3);
NANDC2x1 inst_and_b93_0_0 ( imd_wire93_0_0, A0, A1_inv);
NANDC2x1 inst_and_b93_1_0 ( imd_wire93_1_0, wire93_0_0, wire93_0_1);
NANDC2x1 inst_clockedAND_b92_92 ( imd_YF92, CLK, Y92);
NANDC2x1 inst_and_b92_1_1 ( imd_wire92_1_1, A6, wire92_0_2);
NANDC2x1 inst_and_b92_0_2 ( imd_wire92_0_2, A4, A5_inv);
NANDC2x1 inst_and_b92_2_0 ( imd_Y92, wire92_1_0, wire92_1_1);
NANDC2x1 inst_and_b92_0_1 ( imd_wire92_0_1, A2, A3);
NANDC2x1 inst_and_b92_0_0 ( imd_wire92_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b92_1_0 ( imd_wire92_1_0, wire92_0_0, wire92_0_1);
NANDC2x1 inst_and_b100_1_1 ( imd_wire100_1_1, A6, wire100_0_2);
NANDC2x1 inst_and_b100_0_2 ( imd_wire100_0_2, A4_inv, A5);
NANDC2x1 inst_clockedAND_b91_91 ( imd_YF91, CLK, Y91);
NANDC2x1 inst_and_b91_2_0 ( imd_Y91, wire91_1_0, wire91_1_1);
NANDC2x1 inst_and_b91_0_1 ( imd_wire91_0_1, A2_inv, A3);
NANDC2x1 inst_and_b91_0_0 ( imd_wire91_0_0, A0, A1);
NANDC2x1 inst_and_b91_1_0 ( imd_wire91_1_0, wire91_0_0, wire91_0_1);
NANDC2x1 inst_clockedAND_b90_90 ( imd_YF90, CLK, Y90);
NANDC2x1 inst_and_b90_1_1 ( imd_wire90_1_1, A6, wire90_0_2);
NANDC2x1 inst_and_b90_0_2 ( imd_wire90_0_2, A4, A5_inv);
NANDC2x1 inst_and_b90_2_0 ( imd_Y90, wire90_1_0, wire90_1_1);
NANDC2x1 inst_and_b90_0_1 ( imd_wire90_0_1, A2_inv, A3);
NANDC2x1 inst_and_b90_0_0 ( imd_wire90_0_0, A0_inv, A1);
NANDC2x1 inst_and_b90_1_0 ( imd_wire90_1_0, wire90_0_0, wire90_0_1);
NANDC2x1 inst_clockedAND_b89_89 ( imd_YF89, CLK, Y89);
NANDC2x1 inst_and_b89_1_1 ( imd_wire89_1_1, A6, wire89_0_2);
NANDC2x1 inst_and_b89_0_2 ( imd_wire89_0_2, A4, A5_inv);
NANDC2x1 inst_and_b89_2_0 ( imd_Y89, wire89_1_0, wire89_1_1);
NANDC2x1 inst_and_b89_0_1 ( imd_wire89_0_1, A2_inv, A3);
NANDC2x1 inst_and_b89_0_0 ( imd_wire89_0_0, A0, A1_inv);
NANDC2x1 inst_and_b89_1_0 ( imd_wire89_1_0, wire89_0_0, wire89_0_1);
NANDC2x1 inst_clockedAND_b88_88 ( imd_YF88, CLK, Y88);
NANDC2x1 inst_and_b88_1_1 ( imd_wire88_1_1, A6, wire88_0_2);
NANDC2x1 inst_and_b88_0_2 ( imd_wire88_0_2, A4, A5_inv);
NANDC2x1 inst_and_b88_2_0 ( imd_Y88, wire88_1_0, wire88_1_1);
NANDC2x1 inst_and_b88_0_1 ( imd_wire88_0_1, A2_inv, A3);
NANDC2x1 inst_and_b88_0_0 ( imd_wire88_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b88_1_0 ( imd_wire88_1_0, wire88_0_0, wire88_0_1);
NANDC2x1 inst_clockedAND_b87_87 ( imd_YF87, CLK, Y87);
NANDC2x1 inst_and_b87_1_1 ( imd_wire87_1_1, A6, wire87_0_2);
NANDC2x1 inst_and_b87_0_2 ( imd_wire87_0_2, A4, A5_inv);
NANDC2x1 inst_and_b87_2_0 ( imd_Y87, wire87_1_0, wire87_1_1);
NANDC2x1 inst_and_b87_0_1 ( imd_wire87_0_1, A2, A3_inv);
NANDC2x1 inst_and_b87_0_0 ( imd_wire87_0_0, A0, A1);
NANDC2x1 inst_and_b87_1_0 ( imd_wire87_1_0, wire87_0_0, wire87_0_1);
NANDC2x1 inst_clockedAND_b86_86 ( imd_YF86, CLK, Y86);
NANDC2x1 inst_and_b86_1_1 ( imd_wire86_1_1, A6, wire86_0_2);
NANDC2x1 inst_and_b86_0_2 ( imd_wire86_0_2, A4, A5_inv);
NANDC2x1 inst_and_b86_2_0 ( imd_Y86, wire86_1_0, wire86_1_1);
NANDC2x1 inst_and_b86_0_1 ( imd_wire86_0_1, A2, A3_inv);
NANDC2x1 inst_and_b86_0_0 ( imd_wire86_0_0, A0_inv, A1);
NANDC2x1 inst_and_b86_1_0 ( imd_wire86_1_0, wire86_0_0, wire86_0_1);
NANDC2x1 inst_clockedAND_b85_85 ( imd_YF85, CLK, Y85);
NANDC2x1 inst_and_b85_1_1 ( imd_wire85_1_1, A6, wire85_0_2);
NANDC2x1 inst_and_b85_0_2 ( imd_wire85_0_2, A4, A5_inv);
NANDC2x1 inst_and_b85_2_0 ( imd_Y85, wire85_1_0, wire85_1_1);
NANDC2x1 inst_and_b85_0_1 ( imd_wire85_0_1, A2, A3_inv);
NANDC2x1 inst_and_b85_0_0 ( imd_wire85_0_0, A0, A1_inv);
NANDC2x1 inst_and_b85_1_0 ( imd_wire85_1_0, wire85_0_0, wire85_0_1);
NANDC2x1 inst_clockedAND_b84_84 ( imd_YF84, CLK, Y84);
NANDC2x1 inst_and_b84_1_1 ( imd_wire84_1_1, A6, wire84_0_2);
NANDC2x1 inst_and_b84_0_2 ( imd_wire84_0_2, A4, A5_inv);
NANDC2x1 inst_and_b84_2_0 ( imd_Y84, wire84_1_0, wire84_1_1);
NANDC2x1 inst_and_b84_0_1 ( imd_wire84_0_1, A2, A3_inv);
NANDC2x1 inst_and_b84_0_0 ( imd_wire84_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b84_1_0 ( imd_wire84_1_0, wire84_0_0, wire84_0_1);
NANDC2x1 inst_clockedAND_b83_83 ( imd_YF83, CLK, Y83);
NANDC2x1 inst_and_b83_1_1 ( imd_wire83_1_1, A6, wire83_0_2);
NANDC2x1 inst_and_b83_0_2 ( imd_wire83_0_2, A4, A5_inv);
NANDC2x1 inst_and_b83_2_0 ( imd_Y83, wire83_1_0, wire83_1_1);
NANDC2x1 inst_and_b83_0_1 ( imd_wire83_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b83_0_0 ( imd_wire83_0_0, A0, A1);
NANDC2x1 inst_and_b83_1_0 ( imd_wire83_1_0, wire83_0_0, wire83_0_1);
NANDC2x1 inst_and_b91_1_1 ( imd_wire91_1_1, A6, wire91_0_2);
NANDC2x1 inst_and_b91_0_2 ( imd_wire91_0_2, A4, A5_inv);
NANDC2x1 inst_clockedAND_b82_82 ( imd_YF82, CLK, Y82);
NANDC2x1 inst_and_b82_2_0 ( imd_Y82, wire82_1_0, wire82_1_1);
NANDC2x1 inst_and_b82_0_1 ( imd_wire82_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b82_0_0 ( imd_wire82_0_0, A0_inv, A1);
NANDC2x1 inst_and_b82_1_0 ( imd_wire82_1_0, wire82_0_0, wire82_0_1);
NANDC2x1 inst_clockedAND_b81_81 ( imd_YF81, CLK, Y81);
NANDC2x1 inst_and_b81_1_1 ( imd_wire81_1_1, A6, wire81_0_2);
NANDC2x1 inst_and_b81_0_2 ( imd_wire81_0_2, A4, A5_inv);
NANDC2x1 inst_and_b81_2_0 ( imd_Y81, wire81_1_0, wire81_1_1);
NANDC2x1 inst_and_b81_0_1 ( imd_wire81_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b81_0_0 ( imd_wire81_0_0, A0, A1_inv);
NANDC2x1 inst_and_b81_1_0 ( imd_wire81_1_0, wire81_0_0, wire81_0_1);
NANDC2x1 inst_clockedAND_b80_80 ( imd_YF80, CLK, Y80);
NANDC2x1 inst_and_b80_1_1 ( imd_wire80_1_1, A6, wire80_0_2);
NANDC2x1 inst_and_b80_0_2 ( imd_wire80_0_2, A4, A5_inv);
NANDC2x1 inst_and_b80_2_0 ( imd_Y80, wire80_1_0, wire80_1_1);
NANDC2x1 inst_and_b80_0_1 ( imd_wire80_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b80_0_0 ( imd_wire80_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b80_1_0 ( imd_wire80_1_0, wire80_0_0, wire80_0_1);
NANDC2x1 inst_clockedAND_b79_79 ( imd_YF79, CLK, Y79);
NANDC2x1 inst_and_b79_1_1 ( imd_wire79_1_1, A6, wire79_0_2);
NANDC2x1 inst_and_b79_0_2 ( imd_wire79_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b79_2_0 ( imd_Y79, wire79_1_0, wire79_1_1);
NANDC2x1 inst_and_b79_0_1 ( imd_wire79_0_1, A2, A3);
NANDC2x1 inst_and_b79_0_0 ( imd_wire79_0_0, A0, A1);
NANDC2x1 inst_and_b79_1_0 ( imd_wire79_1_0, wire79_0_0, wire79_0_1);
NANDC2x1 inst_clockedAND_b78_78 ( imd_YF78, CLK, Y78);
NANDC2x1 inst_and_b78_1_1 ( imd_wire78_1_1, A6, wire78_0_2);
NANDC2x1 inst_and_b78_0_2 ( imd_wire78_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b78_2_0 ( imd_Y78, wire78_1_0, wire78_1_1);
NANDC2x1 inst_and_b78_0_1 ( imd_wire78_0_1, A2, A3);
NANDC2x1 inst_and_b78_0_0 ( imd_wire78_0_0, A0_inv, A1);
NANDC2x1 inst_and_b78_1_0 ( imd_wire78_1_0, wire78_0_0, wire78_0_1);
NANDC2x1 inst_clockedAND_b77_77 ( imd_YF77, CLK, Y77);
NANDC2x1 inst_and_b77_1_1 ( imd_wire77_1_1, A6, wire77_0_2);
NANDC2x1 inst_and_b77_0_2 ( imd_wire77_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b77_2_0 ( imd_Y77, wire77_1_0, wire77_1_1);
NANDC2x1 inst_and_b77_0_1 ( imd_wire77_0_1, A2, A3);
NANDC2x1 inst_and_b77_0_0 ( imd_wire77_0_0, A0, A1_inv);
NANDC2x1 inst_and_b77_1_0 ( imd_wire77_1_0, wire77_0_0, wire77_0_1);
NANDC2x1 inst_clockedAND_b76_76 ( imd_YF76, CLK, Y76);
NANDC2x1 inst_and_b76_1_1 ( imd_wire76_1_1, A6, wire76_0_2);
NANDC2x1 inst_and_b76_0_2 ( imd_wire76_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b76_2_0 ( imd_Y76, wire76_1_0, wire76_1_1);
NANDC2x1 inst_and_b76_0_1 ( imd_wire76_0_1, A2, A3);
NANDC2x1 inst_and_b76_0_0 ( imd_wire76_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b76_1_0 ( imd_wire76_1_0, wire76_0_0, wire76_0_1);
NANDC2x1 inst_clockedAND_b75_75 ( imd_YF75, CLK, Y75);
NANDC2x1 inst_and_b75_1_1 ( imd_wire75_1_1, A6, wire75_0_2);
NANDC2x1 inst_and_b75_0_2 ( imd_wire75_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b75_2_0 ( imd_Y75, wire75_1_0, wire75_1_1);
NANDC2x1 inst_and_b75_0_1 ( imd_wire75_0_1, A2_inv, A3);
NANDC2x1 inst_and_b75_0_0 ( imd_wire75_0_0, A0, A1);
NANDC2x1 inst_and_b75_1_0 ( imd_wire75_1_0, wire75_0_0, wire75_0_1);
NANDC2x1 inst_clockedAND_b74_74 ( imd_YF74, CLK, Y74);
NANDC2x1 inst_and_b74_1_1 ( imd_wire74_1_1, A6, wire74_0_2);
NANDC2x1 inst_and_b74_0_2 ( imd_wire74_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b74_2_0 ( imd_Y74, wire74_1_0, wire74_1_1);
NANDC2x1 inst_and_b74_0_1 ( imd_wire74_0_1, A2_inv, A3);
NANDC2x1 inst_and_b74_0_0 ( imd_wire74_0_0, A0_inv, A1);
NANDC2x1 inst_and_b74_1_0 ( imd_wire74_1_0, wire74_0_0, wire74_0_1);
NANDC2x1 inst_and_b82_1_1 ( imd_wire82_1_1, A6, wire82_0_2);
NANDC2x1 inst_and_b82_0_2 ( imd_wire82_0_2, A4, A5_inv);
NANDC2x1 inst_clockedAND_b73_73 ( imd_YF73, CLK, Y73);
NANDC2x1 inst_and_b73_2_0 ( imd_Y73, wire73_1_0, wire73_1_1);
NANDC2x1 inst_and_b73_0_1 ( imd_wire73_0_1, A2_inv, A3);
NANDC2x1 inst_and_b72_0_1 ( imd_wire72_0_1, A2_inv, A3);
NANDC2x1 inst_and_b73_0_0 ( imd_wire73_0_0, A0, A1_inv);
NANDC2x1 inst_and_b73_1_0 ( imd_wire73_1_0, wire73_0_0, wire73_0_1);
NANDC2x1 inst_clockedAND_b72_72 ( imd_YF72, CLK, Y72);
NANDC2x1 inst_and_b72_1_1 ( imd_wire72_1_1, A6, wire72_0_2);
NANDC2x1 inst_and_b72_0_2 ( imd_wire72_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b72_1_0 ( imd_wire72_1_0, wire72_0_0, wire72_0_1);
NANDC2x1 inst_and_b72_0_0 ( imd_wire72_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b72_2_0 ( imd_Y72, wire72_1_0, wire72_1_1);
NANDC2x1 inst_clockedAND_b71_71 ( imd_YF71, CLK, Y71);
NANDC2x1 inst_and_b71_1_1 ( imd_wire71_1_1, A6, wire71_0_2);
NANDC2x1 inst_and_b71_0_2 ( imd_wire71_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b71_2_0 ( imd_Y71, wire71_1_0, wire71_1_1);
NANDC2x1 inst_and_b71_0_1 ( imd_wire71_0_1, A2, A3_inv);
NANDC2x1 inst_and_b71_0_0 ( imd_wire71_0_0, A0, A1);
NANDC2x1 inst_and_b71_1_0 ( imd_wire71_1_0, wire71_0_0, wire71_0_1);
NANDC2x1 inst_clockedAND_b70_70 ( imd_YF70, CLK, Y70);
NANDC2x1 inst_and_b70_1_1 ( imd_wire70_1_1, A6, wire70_0_2);
NANDC2x1 inst_and_b70_0_2 ( imd_wire70_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b70_2_0 ( imd_Y70, wire70_1_0, wire70_1_1);
NANDC2x1 inst_and_b70_0_1 ( imd_wire70_0_1, A2, A3_inv);
NANDC2x1 inst_and_b70_0_0 ( imd_wire70_0_0, A0_inv, A1);
NANDC2x1 inst_and_b70_1_0 ( imd_wire70_1_0, wire70_0_0, wire70_0_1);
NANDC2x1 inst_clockedAND_b69_69 ( imd_YF69, CLK, Y69);
NANDC2x1 inst_and_b69_1_1 ( imd_wire69_1_1, A6, wire69_0_2);
NANDC2x1 inst_and_b69_0_2 ( imd_wire69_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b69_2_0 ( imd_Y69, wire69_1_0, wire69_1_1);
NANDC2x1 inst_and_b69_0_1 ( imd_wire69_0_1, A2, A3_inv);
NANDC2x1 inst_and_b69_0_0 ( imd_wire69_0_0, A0, A1_inv);
NANDC2x1 inst_and_b69_1_0 ( imd_wire69_1_0, wire69_0_0, wire69_0_1);
NANDC2x1 inst_clockedAND_b68_68 ( imd_YF68, CLK, Y68);
NANDC2x1 inst_and_b68_1_1 ( imd_wire68_1_1, A6, wire68_0_2);
NANDC2x1 inst_and_b68_0_2 ( imd_wire68_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b68_2_0 ( imd_Y68, wire68_1_0, wire68_1_1);
NANDC2x1 inst_and_b68_0_1 ( imd_wire68_0_1, A2, A3_inv);
NANDC2x1 inst_and_b68_0_0 ( imd_wire68_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b68_1_0 ( imd_wire68_1_0, wire68_0_0, wire68_0_1);
NANDC2x1 inst_clockedAND_b67_67 ( imd_YF67, CLK, Y67);
NANDC2x1 inst_and_b67_1_1 ( imd_wire67_1_1, A6, wire67_0_2);
NANDC2x1 inst_and_b67_0_2 ( imd_wire67_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b67_2_0 ( imd_Y67, wire67_1_0, wire67_1_1);
NANDC2x1 inst_and_b67_0_1 ( imd_wire67_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b67_0_0 ( imd_wire67_0_0, A0, A1);
NANDC2x1 inst_and_b67_1_0 ( imd_wire67_1_0, wire67_0_0, wire67_0_1);
NANDC2x1 inst_clockedAND_b66_66 ( imd_YF66, CLK, Y66);
NANDC2x1 inst_and_b66_1_1 ( imd_wire66_1_1, A6, wire66_0_2);
NANDC2x1 inst_and_b66_0_2 ( imd_wire66_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b66_2_0 ( imd_Y66, wire66_1_0, wire66_1_1);
NANDC2x1 inst_and_b66_0_1 ( imd_wire66_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b66_0_0 ( imd_wire66_0_0, A0_inv, A1);
NANDC2x1 inst_and_b66_1_0 ( imd_wire66_1_0, wire66_0_0, wire66_0_1);
NANDC2x1 inst_clockedAND_b65_65 ( imd_YF65, CLK, Y65);
NANDC2x1 inst_and_b65_1_1 ( imd_wire65_1_1, A6, wire65_0_2);
NANDC2x1 inst_and_b65_0_2 ( imd_wire65_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b65_2_0 ( imd_Y65, wire65_1_0, wire65_1_1);
NANDC2x1 inst_and_b65_0_1 ( imd_wire65_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b65_0_0 ( imd_wire65_0_0, A0, A1_inv);
NANDC2x1 inst_and_b65_1_0 ( imd_wire65_1_0, wire65_0_0, wire65_0_1);
NANDC2x1 inst_and_b73_1_1 ( imd_wire73_1_1, A6, wire73_0_2);
NANDC2x1 inst_and_b73_0_2 ( imd_wire73_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b64_1_1 ( imd_wire64_1_1, A6, wire64_0_2);
NANDC2x1 inst_and_b64_0_2 ( imd_wire64_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b64_0_1 ( imd_wire64_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b64_0_0 ( imd_wire64_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b64_1_0 ( imd_wire64_1_0, wire64_0_0, wire64_0_1);
NANDC2x1 inst_clockedAND_b63_63 ( imd_YF63, CLK, Y63);
NANDC2x1 inst_and_b63_1_1 ( imd_wire63_1_1, A6_inv, wire63_0_2);
NANDC2x1 inst_and_b63_0_2 ( imd_wire63_0_2, A4, A5);
NANDC2x1 inst_and_b63_2_0 ( imd_Y63, wire63_1_0, wire63_1_1);
NANDC2x1 inst_and_b63_0_1 ( imd_wire63_0_1, A2, A3);
NANDC2x1 inst_and_b63_0_0 ( imd_wire63_0_0, A0, A1);
NANDC2x1 inst_and_b63_1_0 ( imd_wire63_1_0, wire63_0_0, wire63_0_1);
NANDC2x1 inst_clockedAND_b62_62 ( imd_YF62, CLK, Y62);
NANDC2x1 inst_and_b62_1_1 ( imd_wire62_1_1, A6_inv, wire62_0_2);
NANDC2x1 inst_and_b62_0_2 ( imd_wire62_0_2, A4, A5);
NANDC2x1 inst_and_b62_2_0 ( imd_Y62, wire62_1_0, wire62_1_1);
NANDC2x1 inst_and_b62_0_1 ( imd_wire62_0_1, A2, A3);
NANDC2x1 inst_and_b62_0_0 ( imd_wire62_0_0, A0_inv, A1);
NANDC2x1 inst_and_b62_1_0 ( imd_wire62_1_0, wire62_0_0, wire62_0_1);
NANDC2x1 inst_clockedAND_b61_61 ( imd_YF61, CLK, Y61);
NANDC2x1 inst_and_b61_1_1 ( imd_wire61_1_1, A6_inv, wire61_0_2);
NANDC2x1 inst_and_b61_0_2 ( imd_wire61_0_2, A4, A5);
NANDC2x1 inst_and_b61_2_0 ( imd_Y61, wire61_1_0, wire61_1_1);
NANDC2x1 inst_and_b61_0_1 ( imd_wire61_0_1, A2, A3);
NANDC2x1 inst_and_b61_0_0 ( imd_wire61_0_0, A0, A1_inv);
NANDC2x1 inst_and_b61_1_0 ( imd_wire61_1_0, wire61_0_0, wire61_0_1);
NANDC2x1 inst_clockedAND_b60_60 ( imd_YF60, CLK, Y60);
NANDC2x1 inst_and_b60_1_1 ( imd_wire60_1_1, A6_inv, wire60_0_2);
NANDC2x1 inst_and_b60_0_2 ( imd_wire60_0_2, A4, A5);
NANDC2x1 inst_and_b60_2_0 ( imd_Y60, wire60_1_0, wire60_1_1);
NANDC2x1 inst_and_b60_0_1 ( imd_wire60_0_1, A2, A3);
NANDC2x1 inst_and_b60_0_0 ( imd_wire60_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b60_1_0 ( imd_wire60_1_0, wire60_0_0, wire60_0_1);
NANDC2x1 inst_clockedAND_b59_59 ( imd_YF59, CLK, Y59);
NANDC2x1 inst_and_b59_1_1 ( imd_wire59_1_1, A6_inv, wire59_0_2);
NANDC2x1 inst_and_b59_0_2 ( imd_wire59_0_2, A4, A5);
NANDC2x1 inst_and_b59_2_0 ( imd_Y59, wire59_1_0, wire59_1_1);
NANDC2x1 inst_and_b59_0_1 ( imd_wire59_0_1, A2_inv, A3);
NANDC2x1 inst_and_b59_0_0 ( imd_wire59_0_0, A0, A1);
NANDC2x1 inst_and_b59_1_0 ( imd_wire59_1_0, wire59_0_0, wire59_0_1);
NANDC2x1 inst_clockedAND_b58_58 ( imd_YF58, CLK, Y58);
NANDC2x1 inst_and_b58_1_1 ( imd_wire58_1_1, A6_inv, wire58_0_2);
NANDC2x1 inst_and_b58_0_2 ( imd_wire58_0_2, A4, A5);
NANDC2x1 inst_and_b58_2_0 ( imd_Y58, wire58_1_0, wire58_1_1);
NANDC2x1 inst_and_b58_0_1 ( imd_wire58_0_1, A2_inv, A3);
NANDC2x1 inst_and_b58_0_0 ( imd_wire58_0_0, A0_inv, A1);
NANDC2x1 inst_and_b58_1_0 ( imd_wire58_1_0, wire58_0_0, wire58_0_1);
NANDC2x1 inst_clockedAND_b57_57 ( imd_YF57, CLK, Y57);
NANDC2x1 inst_and_b57_1_1 ( imd_wire57_1_1, A6_inv, wire57_0_2);
NANDC2x1 inst_and_b57_0_2 ( imd_wire57_0_2, A4, A5);
NANDC2x1 inst_and_b57_2_0 ( imd_Y57, wire57_1_0, wire57_1_1);
NANDC2x1 inst_and_b57_0_1 ( imd_wire57_0_1, A2_inv, A3);
NANDC2x1 inst_and_b57_0_0 ( imd_wire57_0_0, A0, A1_inv);
NANDC2x1 inst_and_b57_1_0 ( imd_wire57_1_0, wire57_0_0, wire57_0_1);
NANDC2x1 inst_clockedAND_b56_56 ( imd_YF56, CLK, Y56);
NANDC2x1 inst_and_b56_1_1 ( imd_wire56_1_1, A6_inv, wire56_0_2);
NANDC2x1 inst_and_b56_0_2 ( imd_wire56_0_2, A4, A5);
NANDC2x1 inst_and_b56_2_0 ( imd_Y56, wire56_1_0, wire56_1_1);
NANDC2x1 inst_and_b56_0_1 ( imd_wire56_0_1, A2_inv, A3);
NANDC2x1 inst_and_b56_0_0 ( imd_wire56_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b56_1_0 ( imd_wire56_1_0, wire56_0_0, wire56_0_1);
NANDC2x1 inst_clockedAND_b64_64 ( imd_YF64, CLK, Y64);
NANDC2x1 inst_and_b64_2_0 ( imd_Y64, wire64_1_0, wire64_1_1);
NANDC2x1 inst_clockedAND_b55_55 ( imd_YF55, CLK, Y55);
NANDC2x1 inst_and_b55_2_0 ( imd_Y55, wire55_1_0, wire55_1_1);
NANDC2x1 inst_and_b55_0_1 ( imd_wire55_0_1, A2, A3_inv);
NANDC2x1 inst_and_b55_0_0 ( imd_wire55_0_0, A0, A1);
NANDC2x1 inst_and_b55_1_0 ( imd_wire55_1_0, wire55_0_0, wire55_0_1);
NANDC2x1 inst_clockedAND_b54_54 ( imd_YF54, CLK, Y54);
NANDC2x1 inst_and_b54_1_1 ( imd_wire54_1_1, A6_inv, wire54_0_2);
NANDC2x1 inst_and_b54_0_2 ( imd_wire54_0_2, A4, A5);
NANDC2x1 inst_and_b54_2_0 ( imd_Y54, wire54_1_0, wire54_1_1);
NANDC2x1 inst_and_b54_0_1 ( imd_wire54_0_1, A2, A3_inv);
NANDC2x1 inst_and_b54_0_0 ( imd_wire54_0_0, A0_inv, A1);
NANDC2x1 inst_and_b54_1_0 ( imd_wire54_1_0, wire54_0_0, wire54_0_1);
NANDC2x1 inst_clockedAND_b53_53 ( imd_YF53, CLK, Y53);
NANDC2x1 inst_and_b53_1_1 ( imd_wire53_1_1, A6_inv, wire53_0_2);
NANDC2x1 inst_and_b53_0_2 ( imd_wire53_0_2, A4, A5);
NANDC2x1 inst_and_b53_2_0 ( imd_Y53, wire53_1_0, wire53_1_1);
NANDC2x1 inst_and_b53_0_1 ( imd_wire53_0_1, A2, A3_inv);
NANDC2x1 inst_and_b53_0_0 ( imd_wire53_0_0, A0, A1_inv);
NANDC2x1 inst_and_b53_1_0 ( imd_wire53_1_0, wire53_0_0, wire53_0_1);
NANDC2x1 inst_clockedAND_b52_52 ( imd_YF52, CLK, Y52);
NANDC2x1 inst_and_b52_1_1 ( imd_wire52_1_1, A6_inv, wire52_0_2);
NANDC2x1 inst_and_b52_0_2 ( imd_wire52_0_2, A4, A5);
NANDC2x1 inst_and_b52_2_0 ( imd_Y52, wire52_1_0, wire52_1_1);
NANDC2x1 inst_and_b52_0_1 ( imd_wire52_0_1, A2, A3_inv);
NANDC2x1 inst_and_b52_0_0 ( imd_wire52_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b52_1_0 ( imd_wire52_1_0, wire52_0_0, wire52_0_1);
NANDC2x1 inst_clockedAND_b51_51 ( imd_YF51, CLK, Y51);
NANDC2x1 inst_and_b51_1_1 ( imd_wire51_1_1, A6_inv, wire51_0_2);
NANDC2x1 inst_and_b51_0_2 ( imd_wire51_0_2, A4, A5);
NANDC2x1 inst_and_b51_2_0 ( imd_Y51, wire51_1_0, wire51_1_1);
NANDC2x1 inst_and_b51_0_1 ( imd_wire51_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b51_0_0 ( imd_wire51_0_0, A0, A1);
NANDC2x1 inst_and_b51_1_0 ( imd_wire51_1_0, wire51_0_0, wire51_0_1);
NANDC2x1 inst_clockedAND_b50_50 ( imd_YF50, CLK, Y50);
NANDC2x1 inst_and_b50_1_1 ( imd_wire50_1_1, A6_inv, wire50_0_2);
NANDC2x1 inst_and_b50_0_2 ( imd_wire50_0_2, A4, A5);
NANDC2x1 inst_and_b50_2_0 ( imd_Y50, wire50_1_0, wire50_1_1);
NANDC2x1 inst_and_b50_0_1 ( imd_wire50_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b50_0_0 ( imd_wire50_0_0, A0_inv, A1);
NANDC2x1 inst_and_b50_1_0 ( imd_wire50_1_0, wire50_0_0, wire50_0_1);
NANDC2x1 inst_clockedAND_b49_49 ( imd_YF49, CLK, Y49);
NANDC2x1 inst_and_b49_1_1 ( imd_wire49_1_1, A6_inv, wire49_0_2);
NANDC2x1 inst_and_b49_0_2 ( imd_wire49_0_2, A4, A5);
NANDC2x1 inst_and_b49_2_0 ( imd_Y49, wire49_1_0, wire49_1_1);
NANDC2x1 inst_and_b49_0_1 ( imd_wire49_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b49_0_0 ( imd_wire49_0_0, A0, A1_inv);
NANDC2x1 inst_and_b49_1_0 ( imd_wire49_1_0, wire49_0_0, wire49_0_1);
NANDC2x1 inst_clockedAND_b48_48 ( imd_YF48, CLK, Y48);
NANDC2x1 inst_and_b48_1_1 ( imd_wire48_1_1, A6_inv, wire48_0_2);
NANDC2x1 inst_and_b48_0_2 ( imd_wire48_0_2, A4, A5);
NANDC2x1 inst_and_b48_2_0 ( imd_Y48, wire48_1_0, wire48_1_1);
NANDC2x1 inst_and_b48_0_1 ( imd_wire48_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b48_0_0 ( imd_wire48_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b48_1_0 ( imd_wire48_1_0, wire48_0_0, wire48_0_1);
NANDC2x1 inst_clockedAND_b47_47 ( imd_YF47, CLK, Y47);
NANDC2x1 inst_and_b47_1_1 ( imd_wire47_1_1, A6_inv, wire47_0_2);
NANDC2x1 inst_and_b47_0_2 ( imd_wire47_0_2, A4_inv, A5);
NANDC2x1 inst_and_b47_2_0 ( imd_Y47, wire47_1_0, wire47_1_1);
NANDC2x1 inst_and_b47_0_1 ( imd_wire47_0_1, A2, A3);
NANDC2x1 inst_and_b47_0_0 ( imd_wire47_0_0, A0, A1);
NANDC2x1 inst_and_b47_1_0 ( imd_wire47_1_0, wire47_0_0, wire47_0_1);
NANDC2x1 inst_and_b55_1_1 ( imd_wire55_1_1, A6_inv, wire55_0_2);
NANDC2x1 inst_and_b55_0_2 ( imd_wire55_0_2, A4, A5);
NANDC2x1 inst_clockedAND_b46_46 ( imd_YF46, CLK, Y46);
NANDC2x1 inst_and_b46_2_0 ( imd_Y46, wire46_1_0, wire46_1_1);
NANDC2x1 inst_and_b46_0_1 ( imd_wire46_0_1, A2, A3);
NANDC2x1 inst_and_b46_0_0 ( imd_wire46_0_0, A0_inv, A1);
NANDC2x1 inst_and_b46_1_0 ( imd_wire46_1_0, wire46_0_0, wire46_0_1);
NANDC2x1 inst_clockedAND_b45_45 ( imd_YF45, CLK, Y45);
NANDC2x1 inst_and_b45_1_1 ( imd_wire45_1_1, A6_inv, wire45_0_2);
NANDC2x1 inst_and_b45_0_2 ( imd_wire45_0_2, A4_inv, A5);
NANDC2x1 inst_and_b45_2_0 ( imd_Y45, wire45_1_0, wire45_1_1);
NANDC2x1 inst_and_b45_0_1 ( imd_wire45_0_1, A2, A3);
NANDC2x1 inst_and_b45_0_0 ( imd_wire45_0_0, A0, A1_inv);
NANDC2x1 inst_and_b45_1_0 ( imd_wire45_1_0, wire45_0_0, wire45_0_1);
NANDC2x1 inst_clockedAND_b44_44 ( imd_YF44, CLK, Y44);
NANDC2x1 inst_and_b44_1_1 ( imd_wire44_1_1, A6_inv, wire44_0_2);
NANDC2x1 inst_and_b44_0_2 ( imd_wire44_0_2, A4_inv, A5);
NANDC2x1 inst_and_b44_2_0 ( imd_Y44, wire44_1_0, wire44_1_1);
NANDC2x1 inst_and_b44_0_1 ( imd_wire44_0_1, A2, A3);
NANDC2x1 inst_and_b44_0_0 ( imd_wire44_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b44_1_0 ( imd_wire44_1_0, wire44_0_0, wire44_0_1);
NANDC2x1 inst_clockedAND_b43_43 ( imd_YF43, CLK, Y43);
NANDC2x1 inst_and_b43_1_1 ( imd_wire43_1_1, A6_inv, wire43_0_2);
NANDC2x1 inst_and_b43_0_2 ( imd_wire43_0_2, A4_inv, A5);
NANDC2x1 inst_and_b43_2_0 ( imd_Y43, wire43_1_0, wire43_1_1);
NANDC2x1 inst_and_b43_0_1 ( imd_wire43_0_1, A2_inv, A3);
NANDC2x1 inst_and_b43_0_0 ( imd_wire43_0_0, A0, A1);
NANDC2x1 inst_and_b43_1_0 ( imd_wire43_1_0, wire43_0_0, wire43_0_1);
NANDC2x1 inst_clockedAND_b42_42 ( imd_YF42, CLK, Y42);
NANDC2x1 inst_and_b42_1_1 ( imd_wire42_1_1, A6_inv, wire42_0_2);
NANDC2x1 inst_and_b42_0_2 ( imd_wire42_0_2, A4_inv, A5);
NANDC2x1 inst_and_b42_2_0 ( imd_Y42, wire42_1_0, wire42_1_1);
NANDC2x1 inst_and_b42_0_1 ( imd_wire42_0_1, A2_inv, A3);
NANDC2x1 inst_and_b42_0_0 ( imd_wire42_0_0, A0_inv, A1);
NANDC2x1 inst_and_b42_1_0 ( imd_wire42_1_0, wire42_0_0, wire42_0_1);
NANDC2x1 inst_clockedAND_b41_41 ( imd_YF41, CLK, Y41);
NANDC2x1 inst_and_b41_1_1 ( imd_wire41_1_1, A6_inv, wire41_0_2);
NANDC2x1 inst_and_b41_0_2 ( imd_wire41_0_2, A4_inv, A5);
NANDC2x1 inst_and_b41_2_0 ( imd_Y41, wire41_1_0, wire41_1_1);
NANDC2x1 inst_and_b41_0_1 ( imd_wire41_0_1, A2_inv, A3);
NANDC2x1 inst_and_b41_0_0 ( imd_wire41_0_0, A0, A1_inv);
NANDC2x1 inst_and_b41_1_0 ( imd_wire41_1_0, wire41_0_0, wire41_0_1);
NANDC2x1 inst_clockedAND_b40_40 ( imd_YF40, CLK, Y40);
NANDC2x1 inst_and_b40_1_1 ( imd_wire40_1_1, A6_inv, wire40_0_2);
NANDC2x1 inst_and_b40_0_2 ( imd_wire40_0_2, A4_inv, A5);
NANDC2x1 inst_and_b40_2_0 ( imd_Y40, wire40_1_0, wire40_1_1);
NANDC2x1 inst_and_b40_0_1 ( imd_wire40_0_1, A2_inv, A3);
NANDC2x1 inst_and_b40_0_0 ( imd_wire40_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b40_1_0 ( imd_wire40_1_0, wire40_0_0, wire40_0_1);
NANDC2x1 inst_clockedAND_b39_39 ( imd_YF39, CLK, Y39);
NANDC2x1 inst_and_b39_1_1 ( imd_wire39_1_1, A6_inv, wire39_0_2);
NANDC2x1 inst_and_b39_0_2 ( imd_wire39_0_2, A4_inv, A5);
NANDC2x1 inst_and_b39_2_0 ( imd_Y39, wire39_1_0, wire39_1_1);
NANDC2x1 inst_and_b39_0_1 ( imd_wire39_0_1, A2, A3_inv);
NANDC2x1 inst_and_b38_0_1 ( imd_wire38_0_1, A2, A3_inv);
NANDC2x1 inst_and_b39_0_0 ( imd_wire39_0_0, A0, A1);
NANDC2x1 inst_and_b39_1_0 ( imd_wire39_1_0, wire39_0_0, wire39_0_1);
NANDC2x1 inst_clockedAND_b38_38 ( imd_YF38, CLK, Y38);
NANDC2x1 inst_and_b38_1_1 ( imd_wire38_1_1, A6_inv, wire38_0_2);
NANDC2x1 inst_and_b38_0_2 ( imd_wire38_0_2, A4_inv, A5);
NANDC2x1 inst_and_b38_1_0 ( imd_wire38_1_0, wire38_0_0, wire38_0_1);
NANDC2x1 inst_and_b38_0_0 ( imd_wire38_0_0, A0_inv, A1);
NANDC2x1 inst_and_b38_2_0 ( imd_Y38, wire38_1_0, wire38_1_1);
NANDC2x1 inst_and_b46_1_1 ( imd_wire46_1_1, A6_inv, wire46_0_2);
NANDC2x1 inst_and_b46_0_2 ( imd_wire46_0_2, A4_inv, A5);
NANDC2x1 inst_clockedAND_b37_37 ( imd_YF37, CLK, Y37);
NANDC2x1 inst_and_b37_2_0 ( imd_Y37, wire37_1_0, wire37_1_1);
NANDC2x1 inst_and_b37_0_1 ( imd_wire37_0_1, A2, A3_inv);
NANDC2x1 inst_and_b37_0_0 ( imd_wire37_0_0, A0, A1_inv);
NANDC2x1 inst_and_b37_1_0 ( imd_wire37_1_0, wire37_0_0, wire37_0_1);
NANDC2x1 inst_clockedAND_b36_36 ( imd_YF36, CLK, Y36);
NANDC2x1 inst_and_b36_1_1 ( imd_wire36_1_1, A6_inv, wire36_0_2);
NANDC2x1 inst_and_b36_0_2 ( imd_wire36_0_2, A4_inv, A5);
NANDC2x1 inst_and_b36_2_0 ( imd_Y36, wire36_1_0, wire36_1_1);
NANDC2x1 inst_and_b36_0_1 ( imd_wire36_0_1, A2, A3_inv);
NANDC2x1 inst_and_b36_0_0 ( imd_wire36_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b36_1_0 ( imd_wire36_1_0, wire36_0_0, wire36_0_1);
NANDC2x1 inst_clockedAND_b35_35 ( imd_YF35, CLK, Y35);
NANDC2x1 inst_and_b35_1_1 ( imd_wire35_1_1, A6_inv, wire35_0_2);
NANDC2x1 inst_and_b35_0_2 ( imd_wire35_0_2, A4_inv, A5);
NANDC2x1 inst_and_b35_2_0 ( imd_Y35, wire35_1_0, wire35_1_1);
NANDC2x1 inst_and_b35_0_1 ( imd_wire35_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b35_0_0 ( imd_wire35_0_0, A0, A1);
NANDC2x1 inst_and_b35_1_0 ( imd_wire35_1_0, wire35_0_0, wire35_0_1);
NANDC2x1 inst_clockedAND_b34_34 ( imd_YF34, CLK, Y34);
NANDC2x1 inst_and_b34_1_1 ( imd_wire34_1_1, A6_inv, wire34_0_2);
NANDC2x1 inst_and_b34_0_2 ( imd_wire34_0_2, A4_inv, A5);
NANDC2x1 inst_and_b34_2_0 ( imd_Y34, wire34_1_0, wire34_1_1);
NANDC2x1 inst_and_b34_0_1 ( imd_wire34_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b34_0_0 ( imd_wire34_0_0, A0_inv, A1);
NANDC2x1 inst_and_b34_1_0 ( imd_wire34_1_0, wire34_0_0, wire34_0_1);
NANDC2x1 inst_clockedAND_b33_33 ( imd_YF33, CLK, Y33);
NANDC2x1 inst_and_b33_1_1 ( imd_wire33_1_1, A6_inv, wire33_0_2);
NANDC2x1 inst_and_b33_0_2 ( imd_wire33_0_2, A4_inv, A5);
NANDC2x1 inst_and_b33_2_0 ( imd_Y33, wire33_1_0, wire33_1_1);
NANDC2x1 inst_and_b33_0_1 ( imd_wire33_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b33_0_0 ( imd_wire33_0_0, A0, A1_inv);
NANDC2x1 inst_and_b33_1_0 ( imd_wire33_1_0, wire33_0_0, wire33_0_1);
NANDC2x1 inst_and_b32_0_2 ( imd_wire32_0_2, A4_inv, A5);
NANDC2x1 inst_and_b32_1_1 ( imd_wire32_1_1, A6_inv, wire32_0_2);
NANDC2x1 inst_clockedAND_b32_32 ( imd_YF32, CLK, Y32);
NANDC2x1 inst_and_b32_2_0 ( imd_Y32, wire32_1_0, wire32_1_1);
NANDC2x1 inst_and_b32_0_1 ( imd_wire32_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b32_0_0 ( imd_wire32_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b32_1_0 ( imd_wire32_1_0, wire32_0_0, wire32_0_1);
NANDC2x1 inst_clockedAND_b31_31 ( imd_YF31, CLK, Y31);
NANDC2x1 inst_and_b31_1_1 ( imd_wire31_1_1, A6_inv, wire31_0_2);
NANDC2x1 inst_and_b31_0_2 ( imd_wire31_0_2, A4, A5_inv);
NANDC2x1 inst_and_b31_2_0 ( imd_Y31, wire31_1_0, wire31_1_1);
NANDC2x1 inst_and_b31_0_1 ( imd_wire31_0_1, A2, A3);
NANDC2x1 inst_and_b31_0_0 ( imd_wire31_0_0, A0, A1);
NANDC2x1 inst_and_b31_1_0 ( imd_wire31_1_0, wire31_0_0, wire31_0_1);
NANDC2x1 inst_clockedAND_b30_30 ( imd_YF30, CLK, Y30);
NANDC2x1 inst_and_b30_1_1 ( imd_wire30_1_1, A6_inv, wire30_0_2);
NANDC2x1 inst_and_b30_0_2 ( imd_wire30_0_2, A4, A5_inv);
NANDC2x1 inst_and_b30_2_0 ( imd_Y30, wire30_1_0, wire30_1_1);
NANDC2x1 inst_and_b30_0_1 ( imd_wire30_0_1, A2, A3);
NANDC2x1 inst_and_b30_0_0 ( imd_wire30_0_0, A0_inv, A1);
NANDC2x1 inst_and_b30_1_0 ( imd_wire30_1_0, wire30_0_0, wire30_0_1);
NANDC2x1 inst_clockedAND_b29_29 ( imd_YF29, CLK, Y29);
NANDC2x1 inst_and_b29_1_1 ( imd_wire29_1_1, A6_inv, wire29_0_2);
NANDC2x1 inst_and_b29_0_2 ( imd_wire29_0_2, A4, A5_inv);
NANDC2x1 inst_and_b29_2_0 ( imd_Y29, wire29_1_0, wire29_1_1);
NANDC2x1 inst_and_b29_0_1 ( imd_wire29_0_1, A2, A3);
NANDC2x1 inst_and_b29_0_0 ( imd_wire29_0_0, A0, A1_inv);
NANDC2x1 inst_and_b29_1_0 ( imd_wire29_1_0, wire29_0_0, wire29_0_1);
NANDC2x1 inst_and_b37_1_1 ( imd_wire37_1_1, A6_inv, wire37_0_2);
NANDC2x1 inst_and_b37_0_2 ( imd_wire37_0_2, A4_inv, A5);
NANDC2x1 inst_clockedAND_b28_28 ( imd_YF28, CLK, Y28);
NANDC2x1 inst_and_b28_2_0 ( imd_Y28, wire28_1_0, wire28_1_1);
NANDC2x1 inst_and_b28_0_1 ( imd_wire28_0_1, A2, A3);
NANDC2x1 inst_and_b28_0_0 ( imd_wire28_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b28_1_0 ( imd_wire28_1_0, wire28_0_0, wire28_0_1);
NANDC2x1 inst_clockedAND_b27_27 ( imd_YF27, CLK, Y27);
NANDC2x1 inst_and_b27_1_1 ( imd_wire27_1_1, A6_inv, wire27_0_2);
NANDC2x1 inst_and_b27_0_2 ( imd_wire27_0_2, A4, A5_inv);
NANDC2x1 inst_and_b27_2_0 ( imd_Y27, wire27_1_0, wire27_1_1);
NANDC2x1 inst_and_b27_0_1 ( imd_wire27_0_1, A2_inv, A3);
NANDC2x1 inst_and_b27_0_0 ( imd_wire27_0_0, A0, A1);
NANDC2x1 inst_and_b27_1_0 ( imd_wire27_1_0, wire27_0_0, wire27_0_1);
NANDC2x1 inst_clockedAND_b26_26 ( imd_YF26, CLK, Y26);
NANDC2x1 inst_and_b26_1_1 ( imd_wire26_1_1, A6_inv, wire26_0_2);
NANDC2x1 inst_and_b26_0_2 ( imd_wire26_0_2, A4, A5_inv);
NANDC2x1 inst_and_b26_2_0 ( imd_Y26, wire26_1_0, wire26_1_1);
NANDC2x1 inst_and_b26_0_1 ( imd_wire26_0_1, A2_inv, A3);
NANDC2x1 inst_and_b26_0_0 ( imd_wire26_0_0, A0_inv, A1);
NANDC2x1 inst_and_b26_1_0 ( imd_wire26_1_0, wire26_0_0, wire26_0_1);
NANDC2x1 inst_clockedAND_b25_25 ( imd_YF25, CLK, Y25);
NANDC2x1 inst_and_b25_1_1 ( imd_wire25_1_1, A6_inv, wire25_0_2);
NANDC2x1 inst_and_b25_0_2 ( imd_wire25_0_2, A4, A5_inv);
NANDC2x1 inst_and_b25_2_0 ( imd_Y25, wire25_1_0, wire25_1_1);
NANDC2x1 inst_and_b25_0_1 ( imd_wire25_0_1, A2_inv, A3);
NANDC2x1 inst_and_b25_0_0 ( imd_wire25_0_0, A0, A1_inv);
NANDC2x1 inst_and_b25_1_0 ( imd_wire25_1_0, wire25_0_0, wire25_0_1);
NANDC2x1 inst_clockedAND_b24_24 ( imd_YF24, CLK, Y24);
NANDC2x1 inst_and_b24_1_1 ( imd_wire24_1_1, A6_inv, wire24_0_2);
NANDC2x1 inst_and_b24_0_2 ( imd_wire24_0_2, A4, A5_inv);
NANDC2x1 inst_and_b24_2_0 ( imd_Y24, wire24_1_0, wire24_1_1);
NANDC2x1 inst_and_b24_0_1 ( imd_wire24_0_1, A2_inv, A3);
NANDC2x1 inst_and_b24_0_0 ( imd_wire24_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b24_1_0 ( imd_wire24_1_0, wire24_0_0, wire24_0_1);
NANDC2x1 inst_clockedAND_b23_23 ( imd_YF23, CLK, Y23);
NANDC2x1 inst_and_b23_1_1 ( imd_wire23_1_1, A6_inv, wire23_0_2);
NANDC2x1 inst_and_b23_0_2 ( imd_wire23_0_2, A4, A5_inv);
NANDC2x1 inst_and_b23_2_0 ( imd_Y23, wire23_1_0, wire23_1_1);
NANDC2x1 inst_and_b23_0_1 ( imd_wire23_0_1, A2, A3_inv);
NANDC2x1 inst_and_b23_0_0 ( imd_wire23_0_0, A0, A1);
NANDC2x1 inst_and_b23_1_0 ( imd_wire23_1_0, wire23_0_0, wire23_0_1);
NANDC2x1 inst_clockedAND_b22_22 ( imd_YF22, CLK, Y22);
NANDC2x1 inst_and_b22_1_1 ( imd_wire22_1_1, A6_inv, wire22_0_2);
NANDC2x1 inst_and_b22_0_2 ( imd_wire22_0_2, A4, A5_inv);
NANDC2x1 inst_and_b22_2_0 ( imd_Y22, wire22_1_0, wire22_1_1);
NANDC2x1 inst_and_b22_0_1 ( imd_wire22_0_1, A2, A3_inv);
NANDC2x1 inst_and_b22_0_0 ( imd_wire22_0_0, A0_inv, A1);
NANDC2x1 inst_and_b22_1_0 ( imd_wire22_1_0, wire22_0_0, wire22_0_1);
NANDC2x1 inst_clockedAND_b21_21 ( imd_YF21, CLK, Y21);
NANDC2x1 inst_and_b21_1_1 ( imd_wire21_1_1, A6_inv, wire21_0_2);
NANDC2x1 inst_and_b21_0_2 ( imd_wire21_0_2, A4, A5_inv);
NANDC2x1 inst_and_b21_2_0 ( imd_Y21, wire21_1_0, wire21_1_1);
NANDC2x1 inst_and_b21_0_1 ( imd_wire21_0_1, A2, A3_inv);
NANDC2x1 inst_and_b21_0_0 ( imd_wire21_0_0, A0, A1_inv);
NANDC2x1 inst_and_b21_1_0 ( imd_wire21_1_0, wire21_0_0, wire21_0_1);
NANDC2x1 inst_clockedAND_b20_20 ( imd_YF20, CLK, Y20);
NANDC2x1 inst_and_b20_1_1 ( imd_wire20_1_1, A6_inv, wire20_0_2);
NANDC2x1 inst_and_b20_0_2 ( imd_wire20_0_2, A4, A5_inv);
NANDC2x1 inst_and_b20_2_0 ( imd_Y20, wire20_1_0, wire20_1_1);
NANDC2x1 inst_and_b20_0_1 ( imd_wire20_0_1, A2, A3_inv);
NANDC2x1 inst_and_b20_0_0 ( imd_wire20_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b20_1_0 ( imd_wire20_1_0, wire20_0_0, wire20_0_1);
NANDC2x1 inst_and_b28_1_1 ( imd_wire28_1_1, A6_inv, wire28_0_2);
NANDC2x1 inst_and_b28_0_2 ( imd_wire28_0_2, A4, A5_inv);
NANDC2x1 inst_clockedAND_b19_19 ( imd_YF19, CLK, Y19);
NANDC2x1 inst_and_b19_2_0 ( imd_Y19, wire19_1_0, wire19_1_1);
NANDC2x1 inst_and_b19_0_1 ( imd_wire19_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b19_0_0 ( imd_wire19_0_0, A0, A1);
NANDC2x1 inst_and_b19_1_0 ( imd_wire19_1_0, wire19_0_0, wire19_0_1);
NANDC2x1 inst_clockedAND_b18_18 ( imd_YF18, CLK, Y18);
NANDC2x1 inst_and_b18_1_1 ( imd_wire18_1_1, A6_inv, wire18_0_2);
NANDC2x1 inst_and_b18_0_2 ( imd_wire18_0_2, A4, A5_inv);
NANDC2x1 inst_and_b18_2_0 ( imd_Y18, wire18_1_0, wire18_1_1);
NANDC2x1 inst_and_b18_0_1 ( imd_wire18_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b18_0_0 ( imd_wire18_0_0, A0_inv, A1);
NANDC2x1 inst_and_b18_1_0 ( imd_wire18_1_0, wire18_0_0, wire18_0_1);
NANDC2x1 inst_clockedAND_b17_17 ( imd_YF17, CLK, Y17);
NANDC2x1 inst_and_b17_1_1 ( imd_wire17_1_1, A6_inv, wire17_0_2);
NANDC2x1 inst_and_b17_0_2 ( imd_wire17_0_2, A4, A5_inv);
NANDC2x1 inst_and_b17_2_0 ( imd_Y17, wire17_1_0, wire17_1_1);
NANDC2x1 inst_and_b17_0_1 ( imd_wire17_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b17_0_0 ( imd_wire17_0_0, A0, A1_inv);
NANDC2x1 inst_and_b17_1_0 ( imd_wire17_1_0, wire17_0_0, wire17_0_1);
NANDC2x1 inst_and_b16_0_2 ( imd_wire16_0_2, A4, A5_inv);
NANDC2x1 inst_and_b16_1_1 ( imd_wire16_1_1, A6_inv, wire16_0_2);
NANDC2x1 inst_clockedAND_b16_16 ( imd_YF16, CLK, Y16);
NANDC2x1 inst_and_b16_2_0 ( imd_Y16, wire16_1_0, wire16_1_1);
NANDC2x1 inst_and_b16_0_1 ( imd_wire16_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b16_0_0 ( imd_wire16_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b16_1_0 ( imd_wire16_1_0, wire16_0_0, wire16_0_1);
NANDC2x1 inst_clockedAND_b15_15 ( imd_YF15, CLK, Y15);
NANDC2x1 inst_and_b15_1_1 ( imd_wire15_1_1, A6_inv, wire15_0_2);
NANDC2x1 inst_and_b15_0_2 ( imd_wire15_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b15_2_0 ( imd_Y15, wire15_1_0, wire15_1_1);
NANDC2x1 inst_and_b15_0_1 ( imd_wire15_0_1, A2, A3);
NANDC2x1 inst_and_b15_0_0 ( imd_wire15_0_0, A0, A1);
NANDC2x1 inst_and_b15_1_0 ( imd_wire15_1_0, wire15_0_0, wire15_0_1);
NANDC2x1 inst_clockedAND_b14_14 ( imd_YF14, CLK, Y14);
NANDC2x1 inst_and_b14_1_1 ( imd_wire14_1_1, A6_inv, wire14_0_2);
NANDC2x1 inst_and_b14_0_2 ( imd_wire14_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b14_2_0 ( imd_Y14, wire14_1_0, wire14_1_1);
NANDC2x1 inst_and_b14_0_1 ( imd_wire14_0_1, A2, A3);
NANDC2x1 inst_and_b14_0_0 ( imd_wire14_0_0, A0_inv, A1);
NANDC2x1 inst_and_b14_1_0 ( imd_wire14_1_0, wire14_0_0, wire14_0_1);
NANDC2x1 inst_clockedAND_b13_13 ( imd_YF13, CLK, Y13);
NANDC2x1 inst_and_b13_1_1 ( imd_wire13_1_1, A6_inv, wire13_0_2);
NANDC2x1 inst_and_b13_0_2 ( imd_wire13_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b13_2_0 ( imd_Y13, wire13_1_0, wire13_1_1);
NANDC2x1 inst_and_b13_0_1 ( imd_wire13_0_1, A2, A3);
NANDC2x1 inst_and_b13_0_0 ( imd_wire13_0_0, A0, A1_inv);
NANDC2x1 inst_and_b13_1_0 ( imd_wire13_1_0, wire13_0_0, wire13_0_1);
NANDC2x1 inst_clockedAND_b12_12 ( imd_YF12, CLK, Y12);
NANDC2x1 inst_and_b12_1_1 ( imd_wire12_1_1, A6_inv, wire12_0_2);
NANDC2x1 inst_and_b12_0_2 ( imd_wire12_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b12_2_0 ( imd_Y12, wire12_1_0, wire12_1_1);
NANDC2x1 inst_and_b12_0_1 ( imd_wire12_0_1, A2, A3);
NANDC2x1 inst_and_b12_0_0 ( imd_wire12_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b12_1_0 ( imd_wire12_1_0, wire12_0_0, wire12_0_1);
NANDC2x1 inst_clockedAND_b11_11 ( imd_YF11, CLK, Y11);
NANDC2x1 inst_and_b11_1_1 ( imd_wire11_1_1, A6_inv, wire11_0_2);
NANDC2x1 inst_and_b11_0_2 ( imd_wire11_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b11_2_0 ( imd_Y11, wire11_1_0, wire11_1_1);
NANDC2x1 inst_and_b11_0_1 ( imd_wire11_0_1, A2_inv, A3);
NANDC2x1 inst_and_b11_0_0 ( imd_wire11_0_0, A0, A1);
NANDC2x1 inst_and_b11_1_0 ( imd_wire11_1_0, wire11_0_0, wire11_0_1);
NANDC2x1 inst_and_b19_1_1 ( imd_wire19_1_1, A6_inv, wire19_0_2);
NANDC2x1 inst_and_b19_0_2 ( imd_wire19_0_2, A4, A5_inv);
NANDC2x1 inst_clockedAND_b10_10 ( imd_YF10, CLK, Y10);
NANDC2x1 inst_and_b10_2_0 ( imd_Y10, wire10_1_0, wire10_1_1);
NANDC2x1 inst_and_b10_0_1 ( imd_wire10_0_1, A2_inv, A3);
NANDC2x1 inst_and_b10_0_0 ( imd_wire10_0_0, A0_inv, A1);
NANDC2x1 inst_and_b10_1_0 ( imd_wire10_1_0, wire10_0_0, wire10_0_1);
NANDC2x1 inst_clockedAND_b9_9 ( imd_YF9, CLK, Y9);
NANDC2x1 inst_and_b9_1_1 ( imd_wire9_1_1, A6_inv, wire9_0_2);
NANDC2x1 inst_and_b9_0_2 ( imd_wire9_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b9_2_0 ( imd_Y9, wire9_1_0, wire9_1_1);
NANDC2x1 inst_and_b9_0_1 ( imd_wire9_0_1, A2_inv, A3);
NANDC2x1 inst_and_b9_0_0 ( imd_wire9_0_0, A0, A1_inv);
NANDC2x1 inst_and_b9_1_0 ( imd_wire9_1_0, wire9_0_0, wire9_0_1);
NANDC2x1 inst_and_b8_0_1 ( imd_wire8_0_1, A2_inv, A3);
NANDC2x1 inst_and_b8_0_0 ( imd_wire8_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b8_1_0 ( imd_wire8_1_0, wire8_0_0, wire8_0_1);
NANDC2x1 inst_clockedAND_b8_8 ( imd_YF8, CLK, Y8);
NANDC2x1 inst_and_b8_1_1 ( imd_wire8_1_1, A6_inv, wire8_0_2);
NANDC2x1 inst_and_b8_0_2 ( imd_wire8_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b8_2_0 ( imd_Y8, wire8_1_0, wire8_1_1);
NANDC2x1 inst_clockedAND_b7_7 ( imd_YF7, CLK, Y7);
NANDC2x1 inst_and_b7_1_1 ( imd_wire7_1_1, A6_inv, wire7_0_2);
NANDC2x1 inst_and_b7_0_2 ( imd_wire7_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b7_2_0 ( imd_Y7, wire7_1_0, wire7_1_1);
NANDC2x1 inst_and_b7_0_1 ( imd_wire7_0_1, A2, A3_inv);
NANDC2x1 inst_and_b7_0_0 ( imd_wire7_0_0, A0, A1);
NANDC2x1 inst_and_b7_1_0 ( imd_wire7_1_0, wire7_0_0, wire7_0_1);
NANDC2x1 inst_clockedAND_b6_6 ( imd_YF6, CLK, Y6);
NANDC2x1 inst_and_b6_1_1 ( imd_wire6_1_1, A6_inv, wire6_0_2);
NANDC2x1 inst_and_b6_0_2 ( imd_wire6_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b6_2_0 ( imd_Y6, wire6_1_0, wire6_1_1);
NANDC2x1 inst_and_b6_0_1 ( imd_wire6_0_1, A2, A3_inv);
NANDC2x1 inst_and_b6_0_0 ( imd_wire6_0_0, A0_inv, A1);
NANDC2x1 inst_and_b6_1_0 ( imd_wire6_1_0, wire6_0_0, wire6_0_1);
NANDC2x1 inst_clockedAND_b5_5 ( imd_YF5, CLK, Y5);
NANDC2x1 inst_and_b5_1_1 ( imd_wire5_1_1, A6_inv, wire5_0_2);
NANDC2x1 inst_and_b5_0_2 ( imd_wire5_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b5_2_0 ( imd_Y5, wire5_1_0, wire5_1_1);
NANDC2x1 inst_and_b5_0_1 ( imd_wire5_0_1, A2, A3_inv);
NANDC2x1 inst_and_b5_0_0 ( imd_wire5_0_0, A0, A1_inv);
NANDC2x1 inst_and_b5_1_0 ( imd_wire5_1_0, wire5_0_0, wire5_0_1);
NANDC2x1 inst_and_b4_0_1 ( imd_wire4_0_1, A2, A3_inv);
NANDC2x1 inst_and_b4_0_0 ( imd_wire4_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b4_1_0 ( imd_wire4_1_0, wire4_0_0, wire4_0_1);
NANDC2x1 inst_clockedAND_b4_4 ( imd_YF4, CLK, Y4);
NANDC2x1 inst_and_b4_1_1 ( imd_wire4_1_1, A6_inv, wire4_0_2);
NANDC2x1 inst_and_b4_0_2 ( imd_wire4_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b4_2_0 ( imd_Y4, wire4_1_0, wire4_1_1);
NANDC2x1 inst_clockedAND_b3_3 ( imd_YF3, CLK, Y3);
NANDC2x1 inst_and_b3_1_1 ( imd_wire3_1_1, A6_inv, wire3_0_2);
NANDC2x1 inst_and_b3_0_2 ( imd_wire3_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b3_2_0 ( imd_Y3, wire3_1_0, wire3_1_1);
NANDC2x1 inst_and_b3_0_1 ( imd_wire3_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b3_0_0 ( imd_wire3_0_0, A0, A1);
NANDC2x1 inst_and_b3_1_0 ( imd_wire3_1_0, wire3_0_0, wire3_0_1);
NANDC2x1 inst_and_b2_0_0 ( imd_wire2_0_0, A0_inv, A1);
NANDC2x1 inst_and_b2_0_1 ( imd_wire2_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b2_1_0 ( imd_wire2_1_0, wire2_0_0, wire2_0_1);
NANDC2x1 inst_clockedAND_b2_2 ( imd_YF2, CLK, Y2);
NANDC2x1 inst_and_b2_1_1 ( imd_wire2_1_1, A6_inv, wire2_0_2);
NANDC2x1 inst_and_b2_0_2 ( imd_wire2_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b2_2_0 ( imd_Y2, wire2_1_0, wire2_1_1);
NANDC2x1 inst_and_b10_1_1 ( imd_wire10_1_1, A6_inv, wire10_0_2);
NANDC2x1 inst_and_b10_0_2 ( imd_wire10_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b1_0_0 ( imd_wire1_0_0, A0, A1_inv);
NANDC2x1 inst_and_b0_0_0 ( imd_wire0_0_0, A0_inv, A1_inv);
NANDC2x1 inst_clockedAND_b1_1 ( imd_YF1, CLK, Y1);
NANDC2x1 inst_and_b1_1_0 ( imd_wire1_1_0, wire1_0_0, wire1_0_1);
NANDC2x1 inst_and_b1_2_0 ( imd_Y1, wire1_1_0, wire1_1_1);
NANDC2x1 inst_and_b1_0_2 ( imd_wire1_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b0_0_2 ( imd_wire0_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b1_1_1 ( imd_wire1_1_1, A6_inv, wire1_0_2);
NANDC2x1 inst_and_b0_1_1 ( imd_wire0_1_1, A6_inv, wire0_0_2);
NANDC2x1 inst_and_b0_1_0 ( imd_wire0_1_0, wire0_0_0, wire0_0_1);
NANDC2x1 inst_and_b1_0_1 ( imd_wire1_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b0_0_1 ( imd_wire0_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b0_2_0 ( imd_Y0, wire0_1_0, wire0_1_1);
NANDC2x1 inst_clockedAND_b0_0 ( imd_YF0, CLK, Y0);
INVC inst_clockedinv_b127_127 ( YF127, imd_YF127);
INVC inst_inv_b127_2_0 ( Y127, imd_Y127);
INVC inst_inv_b127_1_1 ( wire127_1_1, imd_wire127_1_1);
INVC inst_inv_b127_0_2 ( wire127_0_2, imd_wire127_0_2);
INVC inst_inv_b127_1_0 ( wire127_1_0, imd_wire127_1_0);
INVC inst_inv_b127_0_1 ( wire127_0_1, imd_wire127_0_1);
INVC inst_inv_b127_0_0 ( wire127_0_0, imd_wire127_0_0);
INVC inst_clockedinv_b126_126 ( YF126, imd_YF126);
INVC inst_inv_b126_2_0 ( Y126, imd_Y126);
INVC inst_inv_b126_1_1 ( wire126_1_1, imd_wire126_1_1);
INVC inst_inv_b126_0_2 ( wire126_0_2, imd_wire126_0_2);
INVC inst_inv_b126_1_0 ( wire126_1_0, imd_wire126_1_0);
INVC inst_inv_b126_0_1 ( wire126_0_1, imd_wire126_0_1);
INVC inst_inv_b126_0_0 ( wire126_0_0, imd_wire126_0_0);
INVC inst_clockedinv_b125_125 ( YF125, imd_YF125);
INVC inst_inv_b125_2_0 ( Y125, imd_Y125);
INVC inst_inv_b125_1_1 ( wire125_1_1, imd_wire125_1_1);
INVC inst_inv_b125_0_2 ( wire125_0_2, imd_wire125_0_2);
INVC inst_inv_b125_1_0 ( wire125_1_0, imd_wire125_1_0);
INVC inst_inv_b125_0_1 ( wire125_0_1, imd_wire125_0_1);
INVC inst_inv_b125_0_0 ( wire125_0_0, imd_wire125_0_0);
INVC inst_clockedinv_b124_124 ( YF124, imd_YF124);
INVC inst_inv_b124_2_0 ( Y124, imd_Y124);
INVC inst_inv_b124_1_1 ( wire124_1_1, imd_wire124_1_1);
INVC inst_inv_b124_0_2 ( wire124_0_2, imd_wire124_0_2);
INVC inst_inv_b124_1_0 ( wire124_1_0, imd_wire124_1_0);
INVC inst_inv_b124_0_1 ( wire124_0_1, imd_wire124_0_1);
INVC inst_inv_b124_0_0 ( wire124_0_0, imd_wire124_0_0);
INVC inst_clockedinv_b123_123 ( YF123, imd_YF123);
INVC inst_inv_b123_2_0 ( Y123, imd_Y123);
INVC inst_inv_b123_1_1 ( wire123_1_1, imd_wire123_1_1);
INVC inst_inv_b123_0_2 ( wire123_0_2, imd_wire123_0_2);
INVC inst_inv_b123_1_0 ( wire123_1_0, imd_wire123_1_0);
INVC inst_inv_b123_0_1 ( wire123_0_1, imd_wire123_0_1);
INVC inst_inv_b123_0_0 ( wire123_0_0, imd_wire123_0_0);
INVC inst_clockedinv_b122_122 ( YF122, imd_YF122);
INVC inst_inv_b122_2_0 ( Y122, imd_Y122);
INVC inst_inv_b122_1_1 ( wire122_1_1, imd_wire122_1_1);
INVC inst_inv_b122_0_2 ( wire122_0_2, imd_wire122_0_2);
INVC inst_inv_b122_1_0 ( wire122_1_0, imd_wire122_1_0);
INVC inst_inv_b122_0_1 ( wire122_0_1, imd_wire122_0_1);
INVC inst_inv_b122_0_0 ( wire122_0_0, imd_wire122_0_0);
INVC inst_clockedinv_b121_121 ( YF121, imd_YF121);
INVC inst_inv_b121_2_0 ( Y121, imd_Y121);
INVC inst_inv_b121_1_1 ( wire121_1_1, imd_wire121_1_1);
INVC inst_inv_b121_0_2 ( wire121_0_2, imd_wire121_0_2);
INVC inst_inv_b121_1_0 ( wire121_1_0, imd_wire121_1_0);
INVC inst_inv_b121_0_1 ( wire121_0_1, imd_wire121_0_1);
INVC inst_inv_b121_0_0 ( wire121_0_0, imd_wire121_0_0);
INVC inst_clockedinv_b120_120 ( YF120, imd_YF120);
INVC inst_inv_b120_2_0 ( Y120, imd_Y120);
INVC inst_inv_b120_1_1 ( wire120_1_1, imd_wire120_1_1);
INVC inst_inv_b120_0_2 ( wire120_0_2, imd_wire120_0_2);
INVC inst_inv_b120_1_0 ( wire120_1_0, imd_wire120_1_0);
INVC inst_inv_b120_0_1 ( wire120_0_1, imd_wire120_0_1);
INVC inst_inv_b120_0_0 ( wire120_0_0, imd_wire120_0_0);
INVC inst_clockedinv_b119_119 ( YF119, imd_YF119);
INVC inst_inv_b119_2_0 ( Y119, imd_Y119);
INVC inst_inv_b119_1_1 ( wire119_1_1, imd_wire119_1_1);
INVC inst_inv_b119_0_2 ( wire119_0_2, imd_wire119_0_2);
INVC inst_inv_b119_1_0 ( wire119_1_0, imd_wire119_1_0);
INVC inst_inv_b119_0_1 ( wire119_0_1, imd_wire119_0_1);
INVC inst_inv_b119_0_0 ( wire119_0_0, imd_wire119_0_0);
INVC inst_clockedinv_b118_118 ( YF118, imd_YF118);
INVC inst_inv_b118_2_0 ( Y118, imd_Y118);
INVC inst_inv_b118_1_1 ( wire118_1_1, imd_wire118_1_1);
INVC inst_inv_b118_0_2 ( wire118_0_2, imd_wire118_0_2);
INVC inst_inv_b118_1_0 ( wire118_1_0, imd_wire118_1_0);
INVC inst_inv_b118_0_1 ( wire118_0_1, imd_wire118_0_1);
INVC inst_inv_b118_0_0 ( wire118_0_0, imd_wire118_0_0);
INVC inst_clockedinv_b117_117 ( YF117, imd_YF117);
INVC inst_inv_b117_2_0 ( Y117, imd_Y117);
INVC inst_inv_b117_1_1 ( wire117_1_1, imd_wire117_1_1);
INVC inst_inv_b117_0_2 ( wire117_0_2, imd_wire117_0_2);
INVC inst_inv_b117_1_0 ( wire117_1_0, imd_wire117_1_0);
INVC inst_inv_b117_0_1 ( wire117_0_1, imd_wire117_0_1);
INVC inst_inv_b117_0_0 ( wire117_0_0, imd_wire117_0_0);
INVC inst_clockedinv_b116_116 ( YF116, imd_YF116);
INVC inst_inv_b116_2_0 ( Y116, imd_Y116);
INVC inst_inv_b116_1_1 ( wire116_1_1, imd_wire116_1_1);
INVC inst_inv_b116_0_2 ( wire116_0_2, imd_wire116_0_2);
INVC inst_inv_b116_1_0 ( wire116_1_0, imd_wire116_1_0);
INVC inst_inv_b116_0_1 ( wire116_0_1, imd_wire116_0_1);
INVC inst_inv_b116_0_0 ( wire116_0_0, imd_wire116_0_0);
INVC inst_clockedinv_b115_115 ( YF115, imd_YF115);
INVC inst_inv_b115_2_0 ( Y115, imd_Y115);
INVC inst_inv_b115_1_1 ( wire115_1_1, imd_wire115_1_1);
INVC inst_inv_b115_0_2 ( wire115_0_2, imd_wire115_0_2);
INVC inst_inv_b115_1_0 ( wire115_1_0, imd_wire115_1_0);
INVC inst_inv_b115_0_1 ( wire115_0_1, imd_wire115_0_1);
INVC inst_inv_b115_0_0 ( wire115_0_0, imd_wire115_0_0);
INVC inst_clockedinv_b114_114 ( YF114, imd_YF114);
INVC inst_inv_b114_2_0 ( Y114, imd_Y114);
INVC inst_inv_b114_1_1 ( wire114_1_1, imd_wire114_1_1);
INVC inst_inv_b114_0_2 ( wire114_0_2, imd_wire114_0_2);
INVC inst_inv_b114_1_0 ( wire114_1_0, imd_wire114_1_0);
INVC inst_inv_b114_0_1 ( wire114_0_1, imd_wire114_0_1);
INVC inst_inv_b114_0_0 ( wire114_0_0, imd_wire114_0_0);
INVC inst_clockedinv_b113_113 ( YF113, imd_YF113);
INVC inst_inv_b113_2_0 ( Y113, imd_Y113);
INVC inst_inv_b113_1_1 ( wire113_1_1, imd_wire113_1_1);
INVC inst_inv_b113_0_2 ( wire113_0_2, imd_wire113_0_2);
INVC inst_inv_b113_1_0 ( wire113_1_0, imd_wire113_1_0);
INVC inst_inv_b113_0_1 ( wire113_0_1, imd_wire113_0_1);
INVC inst_inv_b113_0_0 ( wire113_0_0, imd_wire113_0_0);
INVC inst_clockedinv_b112_112 ( YF112, imd_YF112);
INVC inst_inv_b112_2_0 ( Y112, imd_Y112);
INVC inst_inv_b112_1_1 ( wire112_1_1, imd_wire112_1_1);
INVC inst_inv_b112_0_2 ( wire112_0_2, imd_wire112_0_2);
INVC inst_inv_b112_1_0 ( wire112_1_0, imd_wire112_1_0);
INVC inst_inv_b112_0_1 ( wire112_0_1, imd_wire112_0_1);
INVC inst_inv_b112_0_0 ( wire112_0_0, imd_wire112_0_0);
INVC inst_inv_b111_1_0 ( wire111_1_0, imd_wire111_1_0);
INVC inst_inv_b111_0_1 ( wire111_0_1, imd_wire111_0_1);
INVC inst_inv_b111_0_0 ( wire111_0_0, imd_wire111_0_0);
INVC inst_clockedinv_b110_110 ( YF110, imd_YF110);
INVC inst_inv_b110_2_0 ( Y110, imd_Y110);
INVC inst_inv_b110_1_1 ( wire110_1_1, imd_wire110_1_1);
INVC inst_inv_b110_1_0 ( wire110_1_0, imd_wire110_1_0);
INVC inst_inv_b110_0_0 ( wire110_0_0, imd_wire110_0_0);
INVC inst_clockedinv_b111_111 ( YF111, imd_YF111);
INVC inst_inv_b111_2_0 ( Y111, imd_Y111);
INVC inst_inv_b111_0_2 ( wire111_0_2, imd_wire111_0_2);
INVC inst_inv_b111_1_1 ( wire111_1_1, imd_wire111_1_1);
INVC inst_inv_b110_0_2 ( wire110_0_2, imd_wire110_0_2);
INVC inst_inv_b110_0_1 ( wire110_0_1, imd_wire110_0_1);
INVC inst_clockedinv_b109_109 ( YF109, imd_YF109);
INVC inst_inv_b109_2_0 ( Y109, imd_Y109);
INVC inst_inv_b109_1_1 ( wire109_1_1, imd_wire109_1_1);
INVC inst_inv_b109_0_2 ( wire109_0_2, imd_wire109_0_2);
INVC inst_inv_b109_1_0 ( wire109_1_0, imd_wire109_1_0);
INVC inst_inv_b109_0_1 ( wire109_0_1, imd_wire109_0_1);
INVC inst_inv_b109_0_0 ( wire109_0_0, imd_wire109_0_0);
INVC inst_clockedinv_b108_108 ( YF108, imd_YF108);
INVC inst_inv_b108_2_0 ( Y108, imd_Y108);
INVC inst_inv_b108_1_1 ( wire108_1_1, imd_wire108_1_1);
INVC inst_inv_b108_0_2 ( wire108_0_2, imd_wire108_0_2);
INVC inst_inv_b108_1_0 ( wire108_1_0, imd_wire108_1_0);
INVC inst_inv_b108_0_1 ( wire108_0_1, imd_wire108_0_1);
INVC inst_inv_b108_0_0 ( wire108_0_0, imd_wire108_0_0);
INVC inst_clockedinv_b107_107 ( YF107, imd_YF107);
INVC inst_inv_b107_2_0 ( Y107, imd_Y107);
INVC inst_inv_b107_1_1 ( wire107_1_1, imd_wire107_1_1);
INVC inst_inv_b107_0_2 ( wire107_0_2, imd_wire107_0_2);
INVC inst_inv_b107_1_0 ( wire107_1_0, imd_wire107_1_0);
INVC inst_inv_b107_0_1 ( wire107_0_1, imd_wire107_0_1);
INVC inst_inv_b107_0_0 ( wire107_0_0, imd_wire107_0_0);
INVC inst_clockedinv_b106_106 ( YF106, imd_YF106);
INVC inst_inv_b106_2_0 ( Y106, imd_Y106);
INVC inst_inv_b106_1_1 ( wire106_1_1, imd_wire106_1_1);
INVC inst_inv_b106_0_2 ( wire106_0_2, imd_wire106_0_2);
INVC inst_inv_b106_1_0 ( wire106_1_0, imd_wire106_1_0);
INVC inst_inv_b106_0_1 ( wire106_0_1, imd_wire106_0_1);
INVC inst_inv_b106_0_0 ( wire106_0_0, imd_wire106_0_0);
INVC inst_clockedinv_b105_105 ( YF105, imd_YF105);
INVC inst_inv_b105_2_0 ( Y105, imd_Y105);
INVC inst_inv_b105_1_1 ( wire105_1_1, imd_wire105_1_1);
INVC inst_inv_b105_0_2 ( wire105_0_2, imd_wire105_0_2);
INVC inst_inv_b105_1_0 ( wire105_1_0, imd_wire105_1_0);
INVC inst_inv_b105_0_1 ( wire105_0_1, imd_wire105_0_1);
INVC inst_inv_b105_0_0 ( wire105_0_0, imd_wire105_0_0);
INVC inst_clockedinv_b104_104 ( YF104, imd_YF104);
INVC inst_inv_b104_2_0 ( Y104, imd_Y104);
INVC inst_inv_b104_1_1 ( wire104_1_1, imd_wire104_1_1);
INVC inst_inv_b104_0_2 ( wire104_0_2, imd_wire104_0_2);
INVC inst_inv_b104_1_0 ( wire104_1_0, imd_wire104_1_0);
INVC inst_inv_b104_0_1 ( wire104_0_1, imd_wire104_0_1);
INVC inst_inv_b104_0_0 ( wire104_0_0, imd_wire104_0_0);
INVC inst_clockedinv_b103_103 ( YF103, imd_YF103);
INVC inst_inv_b103_2_0 ( Y103, imd_Y103);
INVC inst_inv_b103_1_1 ( wire103_1_1, imd_wire103_1_1);
INVC inst_inv_b103_0_2 ( wire103_0_2, imd_wire103_0_2);
INVC inst_inv_b103_1_0 ( wire103_1_0, imd_wire103_1_0);
INVC inst_inv_b103_0_1 ( wire103_0_1, imd_wire103_0_1);
INVC inst_inv_b103_0_0 ( wire103_0_0, imd_wire103_0_0);
INVC inst_clockedinv_b102_102 ( YF102, imd_YF102);
INVC inst_inv_b102_2_0 ( Y102, imd_Y102);
INVC inst_inv_b102_1_1 ( wire102_1_1, imd_wire102_1_1);
INVC inst_inv_b102_0_2 ( wire102_0_2, imd_wire102_0_2);
INVC inst_inv_b102_1_0 ( wire102_1_0, imd_wire102_1_0);
INVC inst_inv_b102_0_1 ( wire102_0_1, imd_wire102_0_1);
INVC inst_inv_b102_0_0 ( wire102_0_0, imd_wire102_0_0);
INVC inst_clockedinv_b101_101 ( YF101, imd_YF101);
INVC inst_inv_b101_2_0 ( Y101, imd_Y101);
INVC inst_inv_b101_1_1 ( wire101_1_1, imd_wire101_1_1);
INVC inst_inv_b101_0_2 ( wire101_0_2, imd_wire101_0_2);
INVC inst_inv_b101_1_0 ( wire101_1_0, imd_wire101_1_0);
INVC inst_inv_b101_0_1 ( wire101_0_1, imd_wire101_0_1);
INVC inst_inv_b101_0_0 ( wire101_0_0, imd_wire101_0_0);
INVC inst_clockedinv_b100_100 ( YF100, imd_YF100);
INVC inst_inv_b100_2_0 ( Y100, imd_Y100);
INVC inst_inv_b100_1_0 ( wire100_1_0, imd_wire100_1_0);
INVC inst_inv_b100_0_1 ( wire100_0_1, imd_wire100_0_1);
INVC inst_inv_b100_0_0 ( wire100_0_0, imd_wire100_0_0);
INVC inst_clockedinv_b99_99 ( YF99, imd_YF99);
INVC inst_inv_b99_2_0 ( Y99, imd_Y99);
INVC inst_inv_b99_1_1 ( wire99_1_1, imd_wire99_1_1);
INVC inst_inv_b99_0_2 ( wire99_0_2, imd_wire99_0_2);
INVC inst_inv_b99_1_0 ( wire99_1_0, imd_wire99_1_0);
INVC inst_inv_b99_0_1 ( wire99_0_1, imd_wire99_0_1);
INVC inst_inv_b99_0_0 ( wire99_0_0, imd_wire99_0_0);
INVC inst_clockedinv_b98_98 ( YF98, imd_YF98);
INVC inst_inv_b98_2_0 ( Y98, imd_Y98);
INVC inst_inv_b98_1_1 ( wire98_1_1, imd_wire98_1_1);
INVC inst_inv_b98_0_2 ( wire98_0_2, imd_wire98_0_2);
INVC inst_inv_b98_1_0 ( wire98_1_0, imd_wire98_1_0);
INVC inst_inv_b98_0_1 ( wire98_0_1, imd_wire98_0_1);
INVC inst_inv_b98_0_0 ( wire98_0_0, imd_wire98_0_0);
INVC inst_clockedinv_b97_97 ( YF97, imd_YF97);
INVC inst_inv_b97_2_0 ( Y97, imd_Y97);
INVC inst_inv_b97_1_1 ( wire97_1_1, imd_wire97_1_1);
INVC inst_inv_b97_0_2 ( wire97_0_2, imd_wire97_0_2);
INVC inst_inv_b97_1_0 ( wire97_1_0, imd_wire97_1_0);
INVC inst_inv_b97_0_1 ( wire97_0_1, imd_wire97_0_1);
INVC inst_inv_b97_0_0 ( wire97_0_0, imd_wire97_0_0);
INVC inst_clockedinv_b96_96 ( YF96, imd_YF96);
INVC inst_inv_b96_2_0 ( Y96, imd_Y96);
INVC inst_inv_b96_1_1 ( wire96_1_1, imd_wire96_1_1);
INVC inst_inv_b96_0_2 ( wire96_0_2, imd_wire96_0_2);
INVC inst_inv_b96_1_0 ( wire96_1_0, imd_wire96_1_0);
INVC inst_inv_b96_0_1 ( wire96_0_1, imd_wire96_0_1);
INVC inst_inv_b96_0_0 ( wire96_0_0, imd_wire96_0_0);
INVC inst_clockedinv_b95_95 ( YF95, imd_YF95);
INVC inst_inv_b95_2_0 ( Y95, imd_Y95);
INVC inst_inv_b95_1_1 ( wire95_1_1, imd_wire95_1_1);
INVC inst_inv_b95_0_2 ( wire95_0_2, imd_wire95_0_2);
INVC inst_inv_b95_1_0 ( wire95_1_0, imd_wire95_1_0);
INVC inst_inv_b95_0_1 ( wire95_0_1, imd_wire95_0_1);
INVC inst_inv_b95_0_0 ( wire95_0_0, imd_wire95_0_0);
INVC inst_clockedinv_b94_94 ( YF94, imd_YF94);
INVC inst_inv_b94_2_0 ( Y94, imd_Y94);
INVC inst_inv_b94_1_1 ( wire94_1_1, imd_wire94_1_1);
INVC inst_inv_b94_0_2 ( wire94_0_2, imd_wire94_0_2);
INVC inst_inv_b94_1_0 ( wire94_1_0, imd_wire94_1_0);
INVC inst_inv_b94_0_1 ( wire94_0_1, imd_wire94_0_1);
INVC inst_inv_b94_0_0 ( wire94_0_0, imd_wire94_0_0);
INVC inst_clockedinv_b93_93 ( YF93, imd_YF93);
INVC inst_inv_b93_2_0 ( Y93, imd_Y93);
INVC inst_inv_b93_1_1 ( wire93_1_1, imd_wire93_1_1);
INVC inst_inv_b93_0_2 ( wire93_0_2, imd_wire93_0_2);
INVC inst_inv_b93_1_0 ( wire93_1_0, imd_wire93_1_0);
INVC inst_inv_b93_0_1 ( wire93_0_1, imd_wire93_0_1);
INVC inst_inv_b93_0_0 ( wire93_0_0, imd_wire93_0_0);
INVC inst_clockedinv_b92_92 ( YF92, imd_YF92);
INVC inst_inv_b92_2_0 ( Y92, imd_Y92);
INVC inst_inv_b92_1_1 ( wire92_1_1, imd_wire92_1_1);
INVC inst_inv_b92_0_2 ( wire92_0_2, imd_wire92_0_2);
INVC inst_inv_b92_1_0 ( wire92_1_0, imd_wire92_1_0);
INVC inst_inv_b92_0_1 ( wire92_0_1, imd_wire92_0_1);
INVC inst_inv_b92_0_0 ( wire92_0_0, imd_wire92_0_0);
INVC inst_inv_b100_0_2 ( wire100_0_2, imd_wire100_0_2);
INVC inst_inv_b100_1_1 ( wire100_1_1, imd_wire100_1_1);
INVC inst_clockedinv_b91_91 ( YF91, imd_YF91);
INVC inst_inv_b91_2_0 ( Y91, imd_Y91);
INVC inst_inv_b91_1_0 ( wire91_1_0, imd_wire91_1_0);
INVC inst_inv_b91_0_1 ( wire91_0_1, imd_wire91_0_1);
INVC inst_inv_b91_0_0 ( wire91_0_0, imd_wire91_0_0);
INVC inst_clockedinv_b90_90 ( YF90, imd_YF90);
INVC inst_inv_b90_2_0 ( Y90, imd_Y90);
INVC inst_inv_b90_1_1 ( wire90_1_1, imd_wire90_1_1);
INVC inst_inv_b90_0_2 ( wire90_0_2, imd_wire90_0_2);
INVC inst_inv_b90_1_0 ( wire90_1_0, imd_wire90_1_0);
INVC inst_inv_b90_0_1 ( wire90_0_1, imd_wire90_0_1);
INVC inst_inv_b90_0_0 ( wire90_0_0, imd_wire90_0_0);
INVC inst_clockedinv_b89_89 ( YF89, imd_YF89);
INVC inst_inv_b89_2_0 ( Y89, imd_Y89);
INVC inst_inv_b89_1_1 ( wire89_1_1, imd_wire89_1_1);
INVC inst_inv_b89_0_2 ( wire89_0_2, imd_wire89_0_2);
INVC inst_inv_b89_1_0 ( wire89_1_0, imd_wire89_1_0);
INVC inst_inv_b89_0_1 ( wire89_0_1, imd_wire89_0_1);
INVC inst_inv_b89_0_0 ( wire89_0_0, imd_wire89_0_0);
INVC inst_clockedinv_b88_88 ( YF88, imd_YF88);
INVC inst_inv_b88_2_0 ( Y88, imd_Y88);
INVC inst_inv_b88_1_1 ( wire88_1_1, imd_wire88_1_1);
INVC inst_inv_b88_0_2 ( wire88_0_2, imd_wire88_0_2);
INVC inst_inv_b88_1_0 ( wire88_1_0, imd_wire88_1_0);
INVC inst_inv_b88_0_1 ( wire88_0_1, imd_wire88_0_1);
INVC inst_inv_b88_0_0 ( wire88_0_0, imd_wire88_0_0);
INVC inst_clockedinv_b87_87 ( YF87, imd_YF87);
INVC inst_inv_b87_2_0 ( Y87, imd_Y87);
INVC inst_inv_b87_1_1 ( wire87_1_1, imd_wire87_1_1);
INVC inst_inv_b87_0_2 ( wire87_0_2, imd_wire87_0_2);
INVC inst_inv_b87_1_0 ( wire87_1_0, imd_wire87_1_0);
INVC inst_inv_b87_0_1 ( wire87_0_1, imd_wire87_0_1);
INVC inst_inv_b87_0_0 ( wire87_0_0, imd_wire87_0_0);
INVC inst_clockedinv_b86_86 ( YF86, imd_YF86);
INVC inst_inv_b86_2_0 ( Y86, imd_Y86);
INVC inst_inv_b86_1_1 ( wire86_1_1, imd_wire86_1_1);
INVC inst_inv_b86_0_2 ( wire86_0_2, imd_wire86_0_2);
INVC inst_inv_b86_1_0 ( wire86_1_0, imd_wire86_1_0);
INVC inst_inv_b86_0_1 ( wire86_0_1, imd_wire86_0_1);
INVC inst_inv_b86_0_0 ( wire86_0_0, imd_wire86_0_0);
INVC inst_clockedinv_b85_85 ( YF85, imd_YF85);
INVC inst_inv_b85_2_0 ( Y85, imd_Y85);
INVC inst_inv_b85_1_1 ( wire85_1_1, imd_wire85_1_1);
INVC inst_inv_b85_0_2 ( wire85_0_2, imd_wire85_0_2);
INVC inst_inv_b85_1_0 ( wire85_1_0, imd_wire85_1_0);
INVC inst_inv_b85_0_1 ( wire85_0_1, imd_wire85_0_1);
INVC inst_inv_b85_0_0 ( wire85_0_0, imd_wire85_0_0);
INVC inst_clockedinv_b84_84 ( YF84, imd_YF84);
INVC inst_inv_b84_2_0 ( Y84, imd_Y84);
INVC inst_inv_b84_1_1 ( wire84_1_1, imd_wire84_1_1);
INVC inst_inv_b84_0_2 ( wire84_0_2, imd_wire84_0_2);
INVC inst_inv_b84_1_0 ( wire84_1_0, imd_wire84_1_0);
INVC inst_inv_b84_0_1 ( wire84_0_1, imd_wire84_0_1);
INVC inst_inv_b84_0_0 ( wire84_0_0, imd_wire84_0_0);
INVC inst_clockedinv_b83_83 ( YF83, imd_YF83);
INVC inst_inv_b83_2_0 ( Y83, imd_Y83);
INVC inst_inv_b83_1_1 ( wire83_1_1, imd_wire83_1_1);
INVC inst_inv_b83_0_2 ( wire83_0_2, imd_wire83_0_2);
INVC inst_inv_b83_1_0 ( wire83_1_0, imd_wire83_1_0);
INVC inst_inv_b83_0_1 ( wire83_0_1, imd_wire83_0_1);
INVC inst_inv_b83_0_0 ( wire83_0_0, imd_wire83_0_0);
INVC inst_inv_b91_0_2 ( wire91_0_2, imd_wire91_0_2);
INVC inst_inv_b91_1_1 ( wire91_1_1, imd_wire91_1_1);
INVC inst_clockedinv_b82_82 ( YF82, imd_YF82);
INVC inst_inv_b82_2_0 ( Y82, imd_Y82);
INVC inst_inv_b82_1_0 ( wire82_1_0, imd_wire82_1_0);
INVC inst_inv_b82_0_1 ( wire82_0_1, imd_wire82_0_1);
INVC inst_inv_b82_0_0 ( wire82_0_0, imd_wire82_0_0);
INVC inst_clockedinv_b81_81 ( YF81, imd_YF81);
INVC inst_inv_b81_2_0 ( Y81, imd_Y81);
INVC inst_inv_b81_1_1 ( wire81_1_1, imd_wire81_1_1);
INVC inst_inv_b81_0_2 ( wire81_0_2, imd_wire81_0_2);
INVC inst_inv_b81_1_0 ( wire81_1_0, imd_wire81_1_0);
INVC inst_inv_b81_0_1 ( wire81_0_1, imd_wire81_0_1);
INVC inst_inv_b81_0_0 ( wire81_0_0, imd_wire81_0_0);
INVC inst_clockedinv_b80_80 ( YF80, imd_YF80);
INVC inst_inv_b80_2_0 ( Y80, imd_Y80);
INVC inst_inv_b80_1_1 ( wire80_1_1, imd_wire80_1_1);
INVC inst_inv_b80_0_2 ( wire80_0_2, imd_wire80_0_2);
INVC inst_inv_b80_1_0 ( wire80_1_0, imd_wire80_1_0);
INVC inst_inv_b80_0_1 ( wire80_0_1, imd_wire80_0_1);
INVC inst_inv_b80_0_0 ( wire80_0_0, imd_wire80_0_0);
INVC inst_clockedinv_b79_79 ( YF79, imd_YF79);
INVC inst_inv_b79_2_0 ( Y79, imd_Y79);
INVC inst_inv_b79_1_1 ( wire79_1_1, imd_wire79_1_1);
INVC inst_inv_b79_0_2 ( wire79_0_2, imd_wire79_0_2);
INVC inst_inv_b79_1_0 ( wire79_1_0, imd_wire79_1_0);
INVC inst_inv_b79_0_1 ( wire79_0_1, imd_wire79_0_1);
INVC inst_inv_b79_0_0 ( wire79_0_0, imd_wire79_0_0);
INVC inst_clockedinv_b78_78 ( YF78, imd_YF78);
INVC inst_inv_b78_2_0 ( Y78, imd_Y78);
INVC inst_inv_b78_1_1 ( wire78_1_1, imd_wire78_1_1);
INVC inst_inv_b78_0_2 ( wire78_0_2, imd_wire78_0_2);
INVC inst_inv_b78_1_0 ( wire78_1_0, imd_wire78_1_0);
INVC inst_inv_b78_0_1 ( wire78_0_1, imd_wire78_0_1);
INVC inst_inv_b78_0_0 ( wire78_0_0, imd_wire78_0_0);
INVC inst_clockedinv_b77_77 ( YF77, imd_YF77);
INVC inst_inv_b77_2_0 ( Y77, imd_Y77);
INVC inst_inv_b77_1_1 ( wire77_1_1, imd_wire77_1_1);
INVC inst_inv_b77_0_2 ( wire77_0_2, imd_wire77_0_2);
INVC inst_inv_b77_1_0 ( wire77_1_0, imd_wire77_1_0);
INVC inst_inv_b77_0_1 ( wire77_0_1, imd_wire77_0_1);
INVC inst_inv_b77_0_0 ( wire77_0_0, imd_wire77_0_0);
INVC inst_clockedinv_b76_76 ( YF76, imd_YF76);
INVC inst_inv_b76_2_0 ( Y76, imd_Y76);
INVC inst_inv_b76_1_1 ( wire76_1_1, imd_wire76_1_1);
INVC inst_inv_b76_0_2 ( wire76_0_2, imd_wire76_0_2);
INVC inst_inv_b76_1_0 ( wire76_1_0, imd_wire76_1_0);
INVC inst_inv_b76_0_1 ( wire76_0_1, imd_wire76_0_1);
INVC inst_inv_b76_0_0 ( wire76_0_0, imd_wire76_0_0);
INVC inst_clockedinv_b75_75 ( YF75, imd_YF75);
INVC inst_inv_b75_2_0 ( Y75, imd_Y75);
INVC inst_inv_b75_1_1 ( wire75_1_1, imd_wire75_1_1);
INVC inst_inv_b75_0_2 ( wire75_0_2, imd_wire75_0_2);
INVC inst_inv_b75_1_0 ( wire75_1_0, imd_wire75_1_0);
INVC inst_inv_b75_0_1 ( wire75_0_1, imd_wire75_0_1);
INVC inst_inv_b75_0_0 ( wire75_0_0, imd_wire75_0_0);
INVC inst_clockedinv_b74_74 ( YF74, imd_YF74);
INVC inst_inv_b74_2_0 ( Y74, imd_Y74);
INVC inst_inv_b74_1_1 ( wire74_1_1, imd_wire74_1_1);
INVC inst_inv_b74_0_2 ( wire74_0_2, imd_wire74_0_2);
INVC inst_inv_b74_1_0 ( wire74_1_0, imd_wire74_1_0);
INVC inst_inv_b74_0_1 ( wire74_0_1, imd_wire74_0_1);
INVC inst_inv_b74_0_0 ( wire74_0_0, imd_wire74_0_0);
INVC inst_inv_b82_0_2 ( wire82_0_2, imd_wire82_0_2);
INVC inst_inv_b82_1_1 ( wire82_1_1, imd_wire82_1_1);
INVC inst_clockedinv_b73_73 ( YF73, imd_YF73);
INVC inst_inv_b73_2_0 ( Y73, imd_Y73);
INVC inst_inv_b73_1_0 ( wire73_1_0, imd_wire73_1_0);
INVC inst_inv_b73_0_1 ( wire73_0_1, imd_wire73_0_1);
INVC inst_inv_b73_0_0 ( wire73_0_0, imd_wire73_0_0);
INVC inst_clockedinv_b72_72 ( YF72, imd_YF72);
INVC inst_inv_b72_2_0 ( Y72, imd_Y72);
INVC inst_inv_b72_1_1 ( wire72_1_1, imd_wire72_1_1);
INVC inst_inv_b72_0_2 ( wire72_0_2, imd_wire72_0_2);
INVC inst_inv_b72_1_0 ( wire72_1_0, imd_wire72_1_0);
INVC inst_inv_b72_0_0 ( wire72_0_0, imd_wire72_0_0);
INVC inst_inv_b72_0_1 ( wire72_0_1, imd_wire72_0_1);
INVC inst_clockedinv_b71_71 ( YF71, imd_YF71);
INVC inst_inv_b71_2_0 ( Y71, imd_Y71);
INVC inst_inv_b71_1_1 ( wire71_1_1, imd_wire71_1_1);
INVC inst_inv_b71_0_2 ( wire71_0_2, imd_wire71_0_2);
INVC inst_inv_b71_1_0 ( wire71_1_0, imd_wire71_1_0);
INVC inst_inv_b71_0_1 ( wire71_0_1, imd_wire71_0_1);
INVC inst_inv_b71_0_0 ( wire71_0_0, imd_wire71_0_0);
INVC inst_clockedinv_b70_70 ( YF70, imd_YF70);
INVC inst_inv_b70_2_0 ( Y70, imd_Y70);
INVC inst_inv_b70_1_1 ( wire70_1_1, imd_wire70_1_1);
INVC inst_inv_b70_0_2 ( wire70_0_2, imd_wire70_0_2);
INVC inst_inv_b70_1_0 ( wire70_1_0, imd_wire70_1_0);
INVC inst_inv_b70_0_1 ( wire70_0_1, imd_wire70_0_1);
INVC inst_inv_b70_0_0 ( wire70_0_0, imd_wire70_0_0);
INVC inst_clockedinv_b69_69 ( YF69, imd_YF69);
INVC inst_inv_b69_2_0 ( Y69, imd_Y69);
INVC inst_inv_b69_1_1 ( wire69_1_1, imd_wire69_1_1);
INVC inst_inv_b69_0_2 ( wire69_0_2, imd_wire69_0_2);
INVC inst_inv_b69_1_0 ( wire69_1_0, imd_wire69_1_0);
INVC inst_inv_b69_0_1 ( wire69_0_1, imd_wire69_0_1);
INVC inst_inv_b69_0_0 ( wire69_0_0, imd_wire69_0_0);
INVC inst_clockedinv_b68_68 ( YF68, imd_YF68);
INVC inst_inv_b68_2_0 ( Y68, imd_Y68);
INVC inst_inv_b68_1_1 ( wire68_1_1, imd_wire68_1_1);
INVC inst_inv_b68_0_2 ( wire68_0_2, imd_wire68_0_2);
INVC inst_inv_b68_1_0 ( wire68_1_0, imd_wire68_1_0);
INVC inst_inv_b68_0_1 ( wire68_0_1, imd_wire68_0_1);
INVC inst_inv_b68_0_0 ( wire68_0_0, imd_wire68_0_0);
INVC inst_clockedinv_b67_67 ( YF67, imd_YF67);
INVC inst_inv_b67_2_0 ( Y67, imd_Y67);
INVC inst_inv_b67_1_1 ( wire67_1_1, imd_wire67_1_1);
INVC inst_inv_b67_0_2 ( wire67_0_2, imd_wire67_0_2);
INVC inst_inv_b67_1_0 ( wire67_1_0, imd_wire67_1_0);
INVC inst_inv_b67_0_1 ( wire67_0_1, imd_wire67_0_1);
INVC inst_inv_b67_0_0 ( wire67_0_0, imd_wire67_0_0);
INVC inst_clockedinv_b66_66 ( YF66, imd_YF66);
INVC inst_inv_b66_2_0 ( Y66, imd_Y66);
INVC inst_inv_b66_1_1 ( wire66_1_1, imd_wire66_1_1);
INVC inst_inv_b66_0_2 ( wire66_0_2, imd_wire66_0_2);
INVC inst_inv_b66_1_0 ( wire66_1_0, imd_wire66_1_0);
INVC inst_inv_b66_0_1 ( wire66_0_1, imd_wire66_0_1);
INVC inst_inv_b66_0_0 ( wire66_0_0, imd_wire66_0_0);
INVC inst_clockedinv_b65_65 ( YF65, imd_YF65);
INVC inst_inv_b65_2_0 ( Y65, imd_Y65);
INVC inst_inv_b65_1_1 ( wire65_1_1, imd_wire65_1_1);
INVC inst_inv_b65_0_2 ( wire65_0_2, imd_wire65_0_2);
INVC inst_inv_b65_1_0 ( wire65_1_0, imd_wire65_1_0);
INVC inst_inv_b65_0_1 ( wire65_0_1, imd_wire65_0_1);
INVC inst_inv_b65_0_0 ( wire65_0_0, imd_wire65_0_0);
INVC inst_inv_b73_0_2 ( wire73_0_2, imd_wire73_0_2);
INVC inst_inv_b73_1_1 ( wire73_1_1, imd_wire73_1_1);
INVC inst_inv_b64_0_2 ( wire64_0_2, imd_wire64_0_2);
INVC inst_inv_b64_1_1 ( wire64_1_1, imd_wire64_1_1);
INVC inst_inv_b64_1_0 ( wire64_1_0, imd_wire64_1_0);
INVC inst_inv_b64_0_1 ( wire64_0_1, imd_wire64_0_1);
INVC inst_inv_b64_0_0 ( wire64_0_0, imd_wire64_0_0);
INVC inst_clockedinv_b63_63 ( YF63, imd_YF63);
INVC inst_inv_b63_2_0 ( Y63, imd_Y63);
INVC inst_inv_b63_1_1 ( wire63_1_1, imd_wire63_1_1);
INVC inst_inv_b63_0_2 ( wire63_0_2, imd_wire63_0_2);
INVC inst_inv_b63_1_0 ( wire63_1_0, imd_wire63_1_0);
INVC inst_inv_b63_0_1 ( wire63_0_1, imd_wire63_0_1);
INVC inst_inv_b63_0_0 ( wire63_0_0, imd_wire63_0_0);
INVC inst_clockedinv_b62_62 ( YF62, imd_YF62);
INVC inst_inv_b62_2_0 ( Y62, imd_Y62);
INVC inst_inv_b62_1_1 ( wire62_1_1, imd_wire62_1_1);
INVC inst_inv_b62_0_2 ( wire62_0_2, imd_wire62_0_2);
INVC inst_inv_b62_1_0 ( wire62_1_0, imd_wire62_1_0);
INVC inst_inv_b62_0_1 ( wire62_0_1, imd_wire62_0_1);
INVC inst_inv_b62_0_0 ( wire62_0_0, imd_wire62_0_0);
INVC inst_clockedinv_b61_61 ( YF61, imd_YF61);
INVC inst_inv_b61_2_0 ( Y61, imd_Y61);
INVC inst_inv_b61_1_1 ( wire61_1_1, imd_wire61_1_1);
INVC inst_inv_b61_0_2 ( wire61_0_2, imd_wire61_0_2);
INVC inst_inv_b61_1_0 ( wire61_1_0, imd_wire61_1_0);
INVC inst_inv_b61_0_1 ( wire61_0_1, imd_wire61_0_1);
INVC inst_inv_b61_0_0 ( wire61_0_0, imd_wire61_0_0);
INVC inst_clockedinv_b60_60 ( YF60, imd_YF60);
INVC inst_inv_b60_2_0 ( Y60, imd_Y60);
INVC inst_inv_b60_1_1 ( wire60_1_1, imd_wire60_1_1);
INVC inst_inv_b60_0_2 ( wire60_0_2, imd_wire60_0_2);
INVC inst_inv_b60_1_0 ( wire60_1_0, imd_wire60_1_0);
INVC inst_inv_b60_0_1 ( wire60_0_1, imd_wire60_0_1);
INVC inst_inv_b60_0_0 ( wire60_0_0, imd_wire60_0_0);
INVC inst_clockedinv_b59_59 ( YF59, imd_YF59);
INVC inst_inv_b59_2_0 ( Y59, imd_Y59);
INVC inst_inv_b59_1_1 ( wire59_1_1, imd_wire59_1_1);
INVC inst_inv_b59_0_2 ( wire59_0_2, imd_wire59_0_2);
INVC inst_inv_b59_1_0 ( wire59_1_0, imd_wire59_1_0);
INVC inst_inv_b59_0_1 ( wire59_0_1, imd_wire59_0_1);
INVC inst_inv_b59_0_0 ( wire59_0_0, imd_wire59_0_0);
INVC inst_clockedinv_b58_58 ( YF58, imd_YF58);
INVC inst_inv_b58_2_0 ( Y58, imd_Y58);
INVC inst_inv_b58_1_1 ( wire58_1_1, imd_wire58_1_1);
INVC inst_inv_b58_0_2 ( wire58_0_2, imd_wire58_0_2);
INVC inst_inv_b58_1_0 ( wire58_1_0, imd_wire58_1_0);
INVC inst_inv_b58_0_1 ( wire58_0_1, imd_wire58_0_1);
INVC inst_inv_b58_0_0 ( wire58_0_0, imd_wire58_0_0);
INVC inst_clockedinv_b57_57 ( YF57, imd_YF57);
INVC inst_inv_b57_2_0 ( Y57, imd_Y57);
INVC inst_inv_b57_1_1 ( wire57_1_1, imd_wire57_1_1);
INVC inst_inv_b57_0_2 ( wire57_0_2, imd_wire57_0_2);
INVC inst_inv_b57_1_0 ( wire57_1_0, imd_wire57_1_0);
INVC inst_inv_b57_0_1 ( wire57_0_1, imd_wire57_0_1);
INVC inst_inv_b57_0_0 ( wire57_0_0, imd_wire57_0_0);
INVC inst_clockedinv_b56_56 ( YF56, imd_YF56);
INVC inst_inv_b56_2_0 ( Y56, imd_Y56);
INVC inst_inv_b56_1_1 ( wire56_1_1, imd_wire56_1_1);
INVC inst_inv_b56_0_2 ( wire56_0_2, imd_wire56_0_2);
INVC inst_inv_b56_1_0 ( wire56_1_0, imd_wire56_1_0);
INVC inst_inv_b56_0_1 ( wire56_0_1, imd_wire56_0_1);
INVC inst_inv_b56_0_0 ( wire56_0_0, imd_wire56_0_0);
INVC inst_clockedinv_b64_64 ( YF64, imd_YF64);
INVC inst_inv_b64_2_0 ( Y64, imd_Y64);
INVC inst_clockedinv_b55_55 ( YF55, imd_YF55);
INVC inst_inv_b55_2_0 ( Y55, imd_Y55);
INVC inst_inv_b55_1_0 ( wire55_1_0, imd_wire55_1_0);
INVC inst_inv_b55_0_1 ( wire55_0_1, imd_wire55_0_1);
INVC inst_inv_b55_0_0 ( wire55_0_0, imd_wire55_0_0);
INVC inst_clockedinv_b54_54 ( YF54, imd_YF54);
INVC inst_inv_b54_2_0 ( Y54, imd_Y54);
INVC inst_inv_b54_1_1 ( wire54_1_1, imd_wire54_1_1);
INVC inst_inv_b54_0_2 ( wire54_0_2, imd_wire54_0_2);
INVC inst_inv_b54_1_0 ( wire54_1_0, imd_wire54_1_0);
INVC inst_inv_b54_0_1 ( wire54_0_1, imd_wire54_0_1);
INVC inst_inv_b54_0_0 ( wire54_0_0, imd_wire54_0_0);
INVC inst_clockedinv_b53_53 ( YF53, imd_YF53);
INVC inst_inv_b53_2_0 ( Y53, imd_Y53);
INVC inst_inv_b53_1_1 ( wire53_1_1, imd_wire53_1_1);
INVC inst_inv_b53_0_2 ( wire53_0_2, imd_wire53_0_2);
INVC inst_inv_b53_1_0 ( wire53_1_0, imd_wire53_1_0);
INVC inst_inv_b53_0_1 ( wire53_0_1, imd_wire53_0_1);
INVC inst_inv_b53_0_0 ( wire53_0_0, imd_wire53_0_0);
INVC inst_clockedinv_b52_52 ( YF52, imd_YF52);
INVC inst_inv_b52_2_0 ( Y52, imd_Y52);
INVC inst_inv_b52_1_1 ( wire52_1_1, imd_wire52_1_1);
INVC inst_inv_b52_0_2 ( wire52_0_2, imd_wire52_0_2);
INVC inst_inv_b52_1_0 ( wire52_1_0, imd_wire52_1_0);
INVC inst_inv_b52_0_1 ( wire52_0_1, imd_wire52_0_1);
INVC inst_inv_b52_0_0 ( wire52_0_0, imd_wire52_0_0);
INVC inst_clockedinv_b51_51 ( YF51, imd_YF51);
INVC inst_inv_b51_2_0 ( Y51, imd_Y51);
INVC inst_inv_b51_1_1 ( wire51_1_1, imd_wire51_1_1);
INVC inst_inv_b51_0_2 ( wire51_0_2, imd_wire51_0_2);
INVC inst_inv_b51_1_0 ( wire51_1_0, imd_wire51_1_0);
INVC inst_inv_b51_0_1 ( wire51_0_1, imd_wire51_0_1);
INVC inst_inv_b51_0_0 ( wire51_0_0, imd_wire51_0_0);
INVC inst_clockedinv_b50_50 ( YF50, imd_YF50);
INVC inst_inv_b50_2_0 ( Y50, imd_Y50);
INVC inst_inv_b50_1_1 ( wire50_1_1, imd_wire50_1_1);
INVC inst_inv_b50_0_2 ( wire50_0_2, imd_wire50_0_2);
INVC inst_inv_b50_1_0 ( wire50_1_0, imd_wire50_1_0);
INVC inst_inv_b50_0_1 ( wire50_0_1, imd_wire50_0_1);
INVC inst_inv_b50_0_0 ( wire50_0_0, imd_wire50_0_0);
INVC inst_clockedinv_b49_49 ( YF49, imd_YF49);
INVC inst_inv_b49_2_0 ( Y49, imd_Y49);
INVC inst_inv_b49_1_1 ( wire49_1_1, imd_wire49_1_1);
INVC inst_inv_b49_0_2 ( wire49_0_2, imd_wire49_0_2);
INVC inst_inv_b49_1_0 ( wire49_1_0, imd_wire49_1_0);
INVC inst_inv_b49_0_1 ( wire49_0_1, imd_wire49_0_1);
INVC inst_inv_b49_0_0 ( wire49_0_0, imd_wire49_0_0);
INVC inst_clockedinv_b48_48 ( YF48, imd_YF48);
INVC inst_inv_b48_2_0 ( Y48, imd_Y48);
INVC inst_inv_b48_1_1 ( wire48_1_1, imd_wire48_1_1);
INVC inst_inv_b48_0_2 ( wire48_0_2, imd_wire48_0_2);
INVC inst_inv_b48_1_0 ( wire48_1_0, imd_wire48_1_0);
INVC inst_inv_b48_0_1 ( wire48_0_1, imd_wire48_0_1);
INVC inst_inv_b48_0_0 ( wire48_0_0, imd_wire48_0_0);
INVC inst_clockedinv_b47_47 ( YF47, imd_YF47);
INVC inst_inv_b47_2_0 ( Y47, imd_Y47);
INVC inst_inv_b47_1_1 ( wire47_1_1, imd_wire47_1_1);
INVC inst_inv_b47_0_2 ( wire47_0_2, imd_wire47_0_2);
INVC inst_inv_b47_1_0 ( wire47_1_0, imd_wire47_1_0);
INVC inst_inv_b47_0_1 ( wire47_0_1, imd_wire47_0_1);
INVC inst_inv_b47_0_0 ( wire47_0_0, imd_wire47_0_0);
INVC inst_inv_b55_0_2 ( wire55_0_2, imd_wire55_0_2);
INVC inst_inv_b55_1_1 ( wire55_1_1, imd_wire55_1_1);
INVC inst_clockedinv_b46_46 ( YF46, imd_YF46);
INVC inst_inv_b46_2_0 ( Y46, imd_Y46);
INVC inst_inv_b46_1_0 ( wire46_1_0, imd_wire46_1_0);
INVC inst_inv_b46_0_1 ( wire46_0_1, imd_wire46_0_1);
INVC inst_inv_b46_0_0 ( wire46_0_0, imd_wire46_0_0);
INVC inst_clockedinv_b45_45 ( YF45, imd_YF45);
INVC inst_inv_b45_2_0 ( Y45, imd_Y45);
INVC inst_inv_b45_1_1 ( wire45_1_1, imd_wire45_1_1);
INVC inst_inv_b45_0_2 ( wire45_0_2, imd_wire45_0_2);
INVC inst_inv_b45_1_0 ( wire45_1_0, imd_wire45_1_0);
INVC inst_inv_b45_0_1 ( wire45_0_1, imd_wire45_0_1);
INVC inst_inv_b45_0_0 ( wire45_0_0, imd_wire45_0_0);
INVC inst_clockedinv_b44_44 ( YF44, imd_YF44);
INVC inst_inv_b44_2_0 ( Y44, imd_Y44);
INVC inst_inv_b44_1_1 ( wire44_1_1, imd_wire44_1_1);
INVC inst_inv_b44_0_2 ( wire44_0_2, imd_wire44_0_2);
INVC inst_inv_b44_1_0 ( wire44_1_0, imd_wire44_1_0);
INVC inst_inv_b44_0_1 ( wire44_0_1, imd_wire44_0_1);
INVC inst_inv_b44_0_0 ( wire44_0_0, imd_wire44_0_0);
INVC inst_clockedinv_b43_43 ( YF43, imd_YF43);
INVC inst_inv_b43_2_0 ( Y43, imd_Y43);
INVC inst_inv_b43_1_1 ( wire43_1_1, imd_wire43_1_1);
INVC inst_inv_b43_0_2 ( wire43_0_2, imd_wire43_0_2);
INVC inst_inv_b43_1_0 ( wire43_1_0, imd_wire43_1_0);
INVC inst_inv_b43_0_1 ( wire43_0_1, imd_wire43_0_1);
INVC inst_inv_b43_0_0 ( wire43_0_0, imd_wire43_0_0);
INVC inst_clockedinv_b42_42 ( YF42, imd_YF42);
INVC inst_inv_b42_2_0 ( Y42, imd_Y42);
INVC inst_inv_b42_1_1 ( wire42_1_1, imd_wire42_1_1);
INVC inst_inv_b42_0_2 ( wire42_0_2, imd_wire42_0_2);
INVC inst_inv_b42_1_0 ( wire42_1_0, imd_wire42_1_0);
INVC inst_inv_b42_0_1 ( wire42_0_1, imd_wire42_0_1);
INVC inst_inv_b42_0_0 ( wire42_0_0, imd_wire42_0_0);
INVC inst_clockedinv_b41_41 ( YF41, imd_YF41);
INVC inst_inv_b41_2_0 ( Y41, imd_Y41);
INVC inst_inv_b41_1_1 ( wire41_1_1, imd_wire41_1_1);
INVC inst_inv_b41_0_2 ( wire41_0_2, imd_wire41_0_2);
INVC inst_inv_b41_1_0 ( wire41_1_0, imd_wire41_1_0);
INVC inst_inv_b41_0_1 ( wire41_0_1, imd_wire41_0_1);
INVC inst_inv_b41_0_0 ( wire41_0_0, imd_wire41_0_0);
INVC inst_clockedinv_b40_40 ( YF40, imd_YF40);
INVC inst_inv_b40_2_0 ( Y40, imd_Y40);
INVC inst_inv_b40_1_1 ( wire40_1_1, imd_wire40_1_1);
INVC inst_inv_b40_0_2 ( wire40_0_2, imd_wire40_0_2);
INVC inst_inv_b40_1_0 ( wire40_1_0, imd_wire40_1_0);
INVC inst_inv_b40_0_1 ( wire40_0_1, imd_wire40_0_1);
INVC inst_inv_b40_0_0 ( wire40_0_0, imd_wire40_0_0);
INVC inst_clockedinv_b39_39 ( YF39, imd_YF39);
INVC inst_inv_b39_2_0 ( Y39, imd_Y39);
INVC inst_inv_b39_1_1 ( wire39_1_1, imd_wire39_1_1);
INVC inst_inv_b39_0_2 ( wire39_0_2, imd_wire39_0_2);
INVC inst_inv_b39_1_0 ( wire39_1_0, imd_wire39_1_0);
INVC inst_inv_b39_0_1 ( wire39_0_1, imd_wire39_0_1);
INVC inst_inv_b39_0_0 ( wire39_0_0, imd_wire39_0_0);
INVC inst_clockedinv_b38_38 ( YF38, imd_YF38);
INVC inst_inv_b38_2_0 ( Y38, imd_Y38);
INVC inst_inv_b38_1_1 ( wire38_1_1, imd_wire38_1_1);
INVC inst_inv_b38_0_2 ( wire38_0_2, imd_wire38_0_2);
INVC inst_inv_b38_1_0 ( wire38_1_0, imd_wire38_1_0);
INVC inst_inv_b38_0_0 ( wire38_0_0, imd_wire38_0_0);
INVC inst_inv_b38_0_1 ( wire38_0_1, imd_wire38_0_1);
INVC inst_inv_b46_0_2 ( wire46_0_2, imd_wire46_0_2);
INVC inst_inv_b46_1_1 ( wire46_1_1, imd_wire46_1_1);
INVC inst_clockedinv_b37_37 ( YF37, imd_YF37);
INVC inst_inv_b37_2_0 ( Y37, imd_Y37);
INVC inst_inv_b37_1_0 ( wire37_1_0, imd_wire37_1_0);
INVC inst_inv_b37_0_1 ( wire37_0_1, imd_wire37_0_1);
INVC inst_inv_b37_0_0 ( wire37_0_0, imd_wire37_0_0);
INVC inst_clockedinv_b36_36 ( YF36, imd_YF36);
INVC inst_inv_b36_2_0 ( Y36, imd_Y36);
INVC inst_inv_b36_1_1 ( wire36_1_1, imd_wire36_1_1);
INVC inst_inv_b36_0_2 ( wire36_0_2, imd_wire36_0_2);
INVC inst_inv_b36_1_0 ( wire36_1_0, imd_wire36_1_0);
INVC inst_inv_b36_0_1 ( wire36_0_1, imd_wire36_0_1);
INVC inst_inv_b36_0_0 ( wire36_0_0, imd_wire36_0_0);
INVC inst_clockedinv_b35_35 ( YF35, imd_YF35);
INVC inst_inv_b35_2_0 ( Y35, imd_Y35);
INVC inst_inv_b35_1_1 ( wire35_1_1, imd_wire35_1_1);
INVC inst_inv_b35_0_2 ( wire35_0_2, imd_wire35_0_2);
INVC inst_inv_b35_1_0 ( wire35_1_0, imd_wire35_1_0);
INVC inst_inv_b35_0_1 ( wire35_0_1, imd_wire35_0_1);
INVC inst_inv_b35_0_0 ( wire35_0_0, imd_wire35_0_0);
INVC inst_clockedinv_b34_34 ( YF34, imd_YF34);
INVC inst_inv_b34_2_0 ( Y34, imd_Y34);
INVC inst_inv_b34_1_1 ( wire34_1_1, imd_wire34_1_1);
INVC inst_inv_b34_0_2 ( wire34_0_2, imd_wire34_0_2);
INVC inst_inv_b34_1_0 ( wire34_1_0, imd_wire34_1_0);
INVC inst_inv_b34_0_1 ( wire34_0_1, imd_wire34_0_1);
INVC inst_inv_b34_0_0 ( wire34_0_0, imd_wire34_0_0);
INVC inst_clockedinv_b33_33 ( YF33, imd_YF33);
INVC inst_inv_b33_2_0 ( Y33, imd_Y33);
INVC inst_inv_b33_1_1 ( wire33_1_1, imd_wire33_1_1);
INVC inst_inv_b33_0_2 ( wire33_0_2, imd_wire33_0_2);
INVC inst_inv_b33_1_0 ( wire33_1_0, imd_wire33_1_0);
INVC inst_inv_b33_0_1 ( wire33_0_1, imd_wire33_0_1);
INVC inst_inv_b33_0_0 ( wire33_0_0, imd_wire33_0_0);
INVC inst_inv_b32_0_2 ( wire32_0_2, imd_wire32_0_2);
INVC inst_inv_b32_1_1 ( wire32_1_1, imd_wire32_1_1);
INVC inst_inv_b32_2_0 ( Y32, imd_Y32);
INVC inst_clockedinv_b32_32 ( YF32, imd_YF32);
INVC inst_inv_b32_1_0 ( wire32_1_0, imd_wire32_1_0);
INVC inst_inv_b32_0_1 ( wire32_0_1, imd_wire32_0_1);
INVC inst_inv_b32_0_0 ( wire32_0_0, imd_wire32_0_0);
INVC inst_clockedinv_b31_31 ( YF31, imd_YF31);
INVC inst_inv_b31_2_0 ( Y31, imd_Y31);
INVC inst_inv_b31_1_1 ( wire31_1_1, imd_wire31_1_1);
INVC inst_inv_b31_0_2 ( wire31_0_2, imd_wire31_0_2);
INVC inst_inv_b31_1_0 ( wire31_1_0, imd_wire31_1_0);
INVC inst_inv_b31_0_1 ( wire31_0_1, imd_wire31_0_1);
INVC inst_inv_b31_0_0 ( wire31_0_0, imd_wire31_0_0);
INVC inst_clockedinv_b30_30 ( YF30, imd_YF30);
INVC inst_inv_b30_2_0 ( Y30, imd_Y30);
INVC inst_inv_b30_1_1 ( wire30_1_1, imd_wire30_1_1);
INVC inst_inv_b30_0_2 ( wire30_0_2, imd_wire30_0_2);
INVC inst_inv_b30_1_0 ( wire30_1_0, imd_wire30_1_0);
INVC inst_inv_b30_0_1 ( wire30_0_1, imd_wire30_0_1);
INVC inst_inv_b30_0_0 ( wire30_0_0, imd_wire30_0_0);
INVC inst_clockedinv_b29_29 ( YF29, imd_YF29);
INVC inst_inv_b29_2_0 ( Y29, imd_Y29);
INVC inst_inv_b29_1_1 ( wire29_1_1, imd_wire29_1_1);
INVC inst_inv_b29_0_2 ( wire29_0_2, imd_wire29_0_2);
INVC inst_inv_b29_1_0 ( wire29_1_0, imd_wire29_1_0);
INVC inst_inv_b29_0_1 ( wire29_0_1, imd_wire29_0_1);
INVC inst_inv_b29_0_0 ( wire29_0_0, imd_wire29_0_0);
INVC inst_inv_b37_0_2 ( wire37_0_2, imd_wire37_0_2);
INVC inst_inv_b37_1_1 ( wire37_1_1, imd_wire37_1_1);
INVC inst_clockedinv_b28_28 ( YF28, imd_YF28);
INVC inst_inv_b28_2_0 ( Y28, imd_Y28);
INVC inst_inv_b28_1_0 ( wire28_1_0, imd_wire28_1_0);
INVC inst_inv_b28_0_1 ( wire28_0_1, imd_wire28_0_1);
INVC inst_inv_b28_0_0 ( wire28_0_0, imd_wire28_0_0);
INVC inst_clockedinv_b27_27 ( YF27, imd_YF27);
INVC inst_inv_b27_2_0 ( Y27, imd_Y27);
INVC inst_inv_b27_1_1 ( wire27_1_1, imd_wire27_1_1);
INVC inst_inv_b27_0_2 ( wire27_0_2, imd_wire27_0_2);
INVC inst_inv_b27_1_0 ( wire27_1_0, imd_wire27_1_0);
INVC inst_inv_b27_0_1 ( wire27_0_1, imd_wire27_0_1);
INVC inst_inv_b27_0_0 ( wire27_0_0, imd_wire27_0_0);
INVC inst_clockedinv_b26_26 ( YF26, imd_YF26);
INVC inst_inv_b26_2_0 ( Y26, imd_Y26);
INVC inst_inv_b26_1_1 ( wire26_1_1, imd_wire26_1_1);
INVC inst_inv_b26_0_2 ( wire26_0_2, imd_wire26_0_2);
INVC inst_inv_b26_1_0 ( wire26_1_0, imd_wire26_1_0);
INVC inst_inv_b26_0_1 ( wire26_0_1, imd_wire26_0_1);
INVC inst_inv_b26_0_0 ( wire26_0_0, imd_wire26_0_0);
INVC inst_clockedinv_b25_25 ( YF25, imd_YF25);
INVC inst_inv_b25_2_0 ( Y25, imd_Y25);
INVC inst_inv_b25_1_1 ( wire25_1_1, imd_wire25_1_1);
INVC inst_inv_b25_0_2 ( wire25_0_2, imd_wire25_0_2);
INVC inst_inv_b25_1_0 ( wire25_1_0, imd_wire25_1_0);
INVC inst_inv_b25_0_1 ( wire25_0_1, imd_wire25_0_1);
INVC inst_inv_b25_0_0 ( wire25_0_0, imd_wire25_0_0);
INVC inst_clockedinv_b24_24 ( YF24, imd_YF24);
INVC inst_inv_b24_2_0 ( Y24, imd_Y24);
INVC inst_inv_b24_1_1 ( wire24_1_1, imd_wire24_1_1);
INVC inst_inv_b24_0_2 ( wire24_0_2, imd_wire24_0_2);
INVC inst_inv_b24_1_0 ( wire24_1_0, imd_wire24_1_0);
INVC inst_inv_b24_0_1 ( wire24_0_1, imd_wire24_0_1);
INVC inst_inv_b24_0_0 ( wire24_0_0, imd_wire24_0_0);
INVC inst_clockedinv_b23_23 ( YF23, imd_YF23);
INVC inst_inv_b23_2_0 ( Y23, imd_Y23);
INVC inst_inv_b23_1_1 ( wire23_1_1, imd_wire23_1_1);
INVC inst_inv_b23_0_2 ( wire23_0_2, imd_wire23_0_2);
INVC inst_inv_b23_1_0 ( wire23_1_0, imd_wire23_1_0);
INVC inst_inv_b23_0_1 ( wire23_0_1, imd_wire23_0_1);
INVC inst_inv_b23_0_0 ( wire23_0_0, imd_wire23_0_0);
INVC inst_clockedinv_b22_22 ( YF22, imd_YF22);
INVC inst_inv_b22_2_0 ( Y22, imd_Y22);
INVC inst_inv_b22_1_1 ( wire22_1_1, imd_wire22_1_1);
INVC inst_inv_b22_0_2 ( wire22_0_2, imd_wire22_0_2);
INVC inst_inv_b22_1_0 ( wire22_1_0, imd_wire22_1_0);
INVC inst_inv_b22_0_1 ( wire22_0_1, imd_wire22_0_1);
INVC inst_inv_b22_0_0 ( wire22_0_0, imd_wire22_0_0);
INVC inst_clockedinv_b21_21 ( YF21, imd_YF21);
INVC inst_inv_b21_2_0 ( Y21, imd_Y21);
INVC inst_inv_b21_1_1 ( wire21_1_1, imd_wire21_1_1);
INVC inst_inv_b21_0_2 ( wire21_0_2, imd_wire21_0_2);
INVC inst_inv_b21_1_0 ( wire21_1_0, imd_wire21_1_0);
INVC inst_inv_b21_0_1 ( wire21_0_1, imd_wire21_0_1);
INVC inst_inv_b21_0_0 ( wire21_0_0, imd_wire21_0_0);
INVC inst_clockedinv_b20_20 ( YF20, imd_YF20);
INVC inst_inv_b20_2_0 ( Y20, imd_Y20);
INVC inst_inv_b20_1_1 ( wire20_1_1, imd_wire20_1_1);
INVC inst_inv_b20_0_2 ( wire20_0_2, imd_wire20_0_2);
INVC inst_inv_b20_1_0 ( wire20_1_0, imd_wire20_1_0);
INVC inst_inv_b20_0_1 ( wire20_0_1, imd_wire20_0_1);
INVC inst_inv_b20_0_0 ( wire20_0_0, imd_wire20_0_0);
INVC inst_inv_b28_0_2 ( wire28_0_2, imd_wire28_0_2);
INVC inst_inv_b28_1_1 ( wire28_1_1, imd_wire28_1_1);
INVC inst_clockedinv_b19_19 ( YF19, imd_YF19);
INVC inst_inv_b19_2_0 ( Y19, imd_Y19);
INVC inst_inv_b19_1_0 ( wire19_1_0, imd_wire19_1_0);
INVC inst_inv_b19_0_1 ( wire19_0_1, imd_wire19_0_1);
INVC inst_inv_b19_0_0 ( wire19_0_0, imd_wire19_0_0);
INVC inst_clockedinv_b18_18 ( YF18, imd_YF18);
INVC inst_inv_b18_2_0 ( Y18, imd_Y18);
INVC inst_inv_b18_1_1 ( wire18_1_1, imd_wire18_1_1);
INVC inst_inv_b18_0_2 ( wire18_0_2, imd_wire18_0_2);
INVC inst_inv_b18_1_0 ( wire18_1_0, imd_wire18_1_0);
INVC inst_inv_b18_0_1 ( wire18_0_1, imd_wire18_0_1);
INVC inst_inv_b18_0_0 ( wire18_0_0, imd_wire18_0_0);
INVC inst_clockedinv_b17_17 ( YF17, imd_YF17);
INVC inst_inv_b17_2_0 ( Y17, imd_Y17);
INVC inst_inv_b17_1_1 ( wire17_1_1, imd_wire17_1_1);
INVC inst_inv_b17_0_2 ( wire17_0_2, imd_wire17_0_2);
INVC inst_inv_b17_1_0 ( wire17_1_0, imd_wire17_1_0);
INVC inst_inv_b17_0_1 ( wire17_0_1, imd_wire17_0_1);
INVC inst_inv_b17_0_0 ( wire17_0_0, imd_wire17_0_0);
INVC inst_inv_b16_0_2 ( wire16_0_2, imd_wire16_0_2);
INVC inst_inv_b16_1_1 ( wire16_1_1, imd_wire16_1_1);
INVC inst_inv_b16_2_0 ( Y16, imd_Y16);
INVC inst_clockedinv_b16_16 ( YF16, imd_YF16);
INVC inst_inv_b16_1_0 ( wire16_1_0, imd_wire16_1_0);
INVC inst_inv_b16_0_1 ( wire16_0_1, imd_wire16_0_1);
INVC inst_inv_b16_0_0 ( wire16_0_0, imd_wire16_0_0);
INVC inst_clockedinv_b15_15 ( YF15, imd_YF15);
INVC inst_inv_b15_2_0 ( Y15, imd_Y15);
INVC inst_inv_b15_1_1 ( wire15_1_1, imd_wire15_1_1);
INVC inst_inv_b15_0_2 ( wire15_0_2, imd_wire15_0_2);
INVC inst_inv_b15_1_0 ( wire15_1_0, imd_wire15_1_0);
INVC inst_inv_b15_0_1 ( wire15_0_1, imd_wire15_0_1);
INVC inst_inv_b15_0_0 ( wire15_0_0, imd_wire15_0_0);
INVC inst_clockedinv_b14_14 ( YF14, imd_YF14);
INVC inst_inv_b14_2_0 ( Y14, imd_Y14);
INVC inst_inv_b14_1_1 ( wire14_1_1, imd_wire14_1_1);
INVC inst_inv_b14_0_2 ( wire14_0_2, imd_wire14_0_2);
INVC inst_inv_b14_1_0 ( wire14_1_0, imd_wire14_1_0);
INVC inst_inv_b14_0_1 ( wire14_0_1, imd_wire14_0_1);
INVC inst_inv_b14_0_0 ( wire14_0_0, imd_wire14_0_0);
INVC inst_clockedinv_b13_13 ( YF13, imd_YF13);
INVC inst_inv_b13_2_0 ( Y13, imd_Y13);
INVC inst_inv_b13_1_1 ( wire13_1_1, imd_wire13_1_1);
INVC inst_inv_b13_0_2 ( wire13_0_2, imd_wire13_0_2);
INVC inst_inv_b13_1_0 ( wire13_1_0, imd_wire13_1_0);
INVC inst_inv_b13_0_1 ( wire13_0_1, imd_wire13_0_1);
INVC inst_inv_b13_0_0 ( wire13_0_0, imd_wire13_0_0);
INVC inst_clockedinv_b12_12 ( YF12, imd_YF12);
INVC inst_inv_b12_2_0 ( Y12, imd_Y12);
INVC inst_inv_b12_1_1 ( wire12_1_1, imd_wire12_1_1);
INVC inst_inv_b12_0_2 ( wire12_0_2, imd_wire12_0_2);
INVC inst_inv_b12_1_0 ( wire12_1_0, imd_wire12_1_0);
INVC inst_inv_b12_0_1 ( wire12_0_1, imd_wire12_0_1);
INVC inst_inv_b12_0_0 ( wire12_0_0, imd_wire12_0_0);
INVC inst_clockedinv_b11_11 ( YF11, imd_YF11);
INVC inst_inv_b11_2_0 ( Y11, imd_Y11);
INVC inst_inv_b11_1_1 ( wire11_1_1, imd_wire11_1_1);
INVC inst_inv_b11_0_2 ( wire11_0_2, imd_wire11_0_2);
INVC inst_inv_b11_1_0 ( wire11_1_0, imd_wire11_1_0);
INVC inst_inv_b11_0_1 ( wire11_0_1, imd_wire11_0_1);
INVC inst_inv_b11_0_0 ( wire11_0_0, imd_wire11_0_0);
INVC inst_inv_b19_0_2 ( wire19_0_2, imd_wire19_0_2);
INVC inst_inv_b19_1_1 ( wire19_1_1, imd_wire19_1_1);
INVC inst_clockedinv_b10_10 ( YF10, imd_YF10);
INVC inst_inv_b10_2_0 ( Y10, imd_Y10);
INVC inst_inv_b10_1_0 ( wire10_1_0, imd_wire10_1_0);
INVC inst_inv_b10_0_1 ( wire10_0_1, imd_wire10_0_1);
INVC inst_inv_b10_0_0 ( wire10_0_0, imd_wire10_0_0);
INVC inst_clockedinv_b9_9 ( YF9, imd_YF9);
INVC inst_inv_b9_2_0 ( Y9, imd_Y9);
INVC inst_inv_b9_1_1 ( wire9_1_1, imd_wire9_1_1);
INVC inst_inv_b9_0_2 ( wire9_0_2, imd_wire9_0_2);
INVC inst_inv_b9_1_0 ( wire9_1_0, imd_wire9_1_0);
INVC inst_inv_b9_0_1 ( wire9_0_1, imd_wire9_0_1);
INVC inst_inv_b9_0_0 ( wire9_0_0, imd_wire9_0_0);
INVC inst_inv_b8_0_1 ( wire8_0_1, imd_wire8_0_1);
INVC inst_inv_b8_1_0 ( wire8_1_0, imd_wire8_1_0);
INVC inst_inv_b8_0_0 ( wire8_0_0, imd_wire8_0_0);
INVC inst_inv_b8_2_0 ( Y8, imd_Y8);
INVC inst_clockedinv_b8_8 ( YF8, imd_YF8);
INVC inst_inv_b8_1_1 ( wire8_1_1, imd_wire8_1_1);
INVC inst_inv_b8_0_2 ( wire8_0_2, imd_wire8_0_2);
INVC inst_clockedinv_b7_7 ( YF7, imd_YF7);
INVC inst_inv_b7_2_0 ( Y7, imd_Y7);
INVC inst_inv_b7_1_1 ( wire7_1_1, imd_wire7_1_1);
INVC inst_inv_b7_0_2 ( wire7_0_2, imd_wire7_0_2);
INVC inst_inv_b7_1_0 ( wire7_1_0, imd_wire7_1_0);
INVC inst_inv_b7_0_1 ( wire7_0_1, imd_wire7_0_1);
INVC inst_inv_b7_0_0 ( wire7_0_0, imd_wire7_0_0);
INVC inst_clockedinv_b6_6 ( YF6, imd_YF6);
INVC inst_inv_b6_2_0 ( Y6, imd_Y6);
INVC inst_inv_b6_1_1 ( wire6_1_1, imd_wire6_1_1);
INVC inst_inv_b6_0_2 ( wire6_0_2, imd_wire6_0_2);
INVC inst_inv_b6_1_0 ( wire6_1_0, imd_wire6_1_0);
INVC inst_inv_b6_0_1 ( wire6_0_1, imd_wire6_0_1);
INVC inst_inv_b6_0_0 ( wire6_0_0, imd_wire6_0_0);
INVC inst_clockedinv_b5_5 ( YF5, imd_YF5);
INVC inst_inv_b5_2_0 ( Y5, imd_Y5);
INVC inst_inv_b5_1_1 ( wire5_1_1, imd_wire5_1_1);
INVC inst_inv_b5_0_2 ( wire5_0_2, imd_wire5_0_2);
INVC inst_inv_b5_1_0 ( wire5_1_0, imd_wire5_1_0);
INVC inst_inv_b5_0_1 ( wire5_0_1, imd_wire5_0_1);
INVC inst_inv_b5_0_0 ( wire5_0_0, imd_wire5_0_0);
INVC inst_inv_b4_0_1 ( wire4_0_1, imd_wire4_0_1);
INVC inst_inv_b4_1_0 ( wire4_1_0, imd_wire4_1_0);
INVC inst_inv_b4_0_0 ( wire4_0_0, imd_wire4_0_0);
INVC inst_inv_b4_2_0 ( Y4, imd_Y4);
INVC inst_clockedinv_b4_4 ( YF4, imd_YF4);
INVC inst_inv_b4_1_1 ( wire4_1_1, imd_wire4_1_1);
INVC inst_inv_b4_0_2 ( wire4_0_2, imd_wire4_0_2);
INVC inst_clockedinv_b3_3 ( YF3, imd_YF3);
INVC inst_inv_b3_2_0 ( Y3, imd_Y3);
INVC inst_inv_b3_1_1 ( wire3_1_1, imd_wire3_1_1);
INVC inst_inv_b3_0_2 ( wire3_0_2, imd_wire3_0_2);
INVC inst_inv_b3_1_0 ( wire3_1_0, imd_wire3_1_0);
INVC inst_inv_b3_0_1 ( wire3_0_1, imd_wire3_0_1);
INVC inst_inv_b3_0_0 ( wire3_0_0, imd_wire3_0_0);
INVC inst_inv_b2_0_0 ( wire2_0_0, imd_wire2_0_0);
INVC inst_inv_b2_1_0 ( wire2_1_0, imd_wire2_1_0);
INVC inst_inv_b2_0_1 ( wire2_0_1, imd_wire2_0_1);
INVC inst_inv_b2_2_0 ( Y2, imd_Y2);
INVC inst_clockedinv_b2_2 ( YF2, imd_YF2);
INVC inst_inv_b2_1_1 ( wire2_1_1, imd_wire2_1_1);
INVC inst_inv_b2_0_2 ( wire2_0_2, imd_wire2_0_2);
INVC inst_inv_b10_0_2 ( wire10_0_2, imd_wire10_0_2);
INVC inst_inv_b10_1_1 ( wire10_1_1, imd_wire10_1_1);
INVC inst_inv_b1_0_0 ( wire1_0_0, imd_wire1_0_0);
INVC inst_inv_b0_0_0 ( wire0_0_0, imd_wire0_0_0);
INVC inst_clockedinv_b1_1 ( YF1, imd_YF1);
INVC inst_inv_b1_2_0 ( Y1, imd_Y1);
INVC inst_inv_b1_1_1 ( wire1_1_1, imd_wire1_1_1);
INVC inst_inv_b1_1_0 ( wire1_1_0, imd_wire1_1_0);
INVC inst_inv_b1_0_1 ( wire1_0_1, imd_wire1_0_1);
INVC inst_inv_b1_0_2 ( wire1_0_2, imd_wire1_0_2);
INVC inst_inv_b0_0_2 ( wire0_0_2, imd_wire0_0_2);
INVC inst_inv_b0_1_1 ( wire0_1_1, imd_wire0_1_1);
INVC inst_inv_b0_0_1 ( wire0_0_1, imd_wire0_0_1);
INVC inst_inv_b0_1_0 ( wire0_1_0, imd_wire0_1_0);
INVC inst_inv_b0_2_0 ( Y0, imd_Y0);
INVC inst_clockedinv_b0_0 ( YF0, imd_YF0);

endmodule
// Library - sram_compiled_2kb_r128_c128_w8, Cell -
//sram_compiled_array, View - schematic
// LAST TIME SAVED: Apr 20 20:07:32 2021
// NETLIST TIME: Apr 21 18:57:14 2021
`timescale 1ns / 1ps 

module sram_compiled_array_2kb ( addr0, addr1, addr2, addr3, addr4, addr5,
     addr6, addr7, addr8, addr9, addr10, din0, din1, din2, din3, din4,
     din5, din6, din7, dout0, dout1, dout2, dout3, dout4, dout5, dout6,
     dout7, clk, write_en, sense_en );

output  dout0, dout1, dout2, dout3, dout4, dout5, dout6, dout7;

input  addr0, addr1, addr2, addr3, addr4, addr5, addr6, addr7, addr8,
     addr9, addr10, clk, din0, din1, din2, din3, din4, din5, din6,
     din7, sense_en, write_en;


specify 
    specparam CDS_LIBNAME  = "sram_compiled_2kb_r128_c128_w8";
    specparam CDS_CELLNAME = "sram_compiled_array";
    specparam CDS_VIEWNAME = "schematic";
endspecify

sram_cell_6t_3 inst_cell_127_127 ( BL127, BLN127, WL127);
sram_cell_6t_3 inst_cell_127_126 ( BL126, BLN126, WL127);
sram_cell_6t_3 inst_cell_127_125 ( BL125, BLN125, WL127);
sram_cell_6t_3 inst_cell_127_124 ( BL124, BLN124, WL127);
sram_cell_6t_3 inst_cell_127_123 ( BL123, BLN123, WL127);
sram_cell_6t_3 inst_cell_127_122 ( BL122, BLN122, WL127);
sram_cell_6t_3 inst_cell_127_121 ( BL121, BLN121, WL127);
sram_cell_6t_3 inst_cell_127_120 ( BL120, BLN120, WL127);
sram_cell_6t_3 inst_cell_127_119 ( BL119, BLN119, WL127);
sram_cell_6t_3 inst_cell_127_118 ( BL118, BLN118, WL127);
sram_cell_6t_3 inst_cell_127_117 ( BL117, BLN117, WL127);
sram_cell_6t_3 inst_cell_127_116 ( BL116, BLN116, WL127);
sram_cell_6t_3 inst_cell_127_115 ( BL115, BLN115, WL127);
sram_cell_6t_3 inst_cell_127_114 ( BL114, BLN114, WL127);
sram_cell_6t_3 inst_cell_127_113 ( BL113, BLN113, WL127);
sram_cell_6t_3 inst_cell_127_112 ( BL112, BLN112, WL127);
sram_cell_6t_3 inst_cell_127_111 ( BL111, BLN111, WL127);
sram_cell_6t_3 inst_cell_127_110 ( BL110, BLN110, WL127);
sram_cell_6t_3 inst_cell_127_79 ( BL79, BLN79, WL127);
sram_cell_6t_3 inst_cell_127_78 ( BL78, BLN78, WL127);
sram_cell_6t_3 inst_cell_127_77 ( BL77, BLN77, WL127);
sram_cell_6t_3 inst_cell_127_76 ( BL76, BLN76, WL127);
sram_cell_6t_3 inst_cell_127_75 ( BL75, BLN75, WL127);
sram_cell_6t_3 inst_cell_127_74 ( BL74, BLN74, WL127);
sram_cell_6t_3 inst_cell_127_73 ( BL73, BLN73, WL127);
sram_cell_6t_3 inst_cell_127_72 ( BL72, BLN72, WL127);
sram_cell_6t_3 inst_cell_127_71 ( BL71, BLN71, WL127);
sram_cell_6t_3 inst_cell_127_70 ( BL70, BLN70, WL127);
sram_cell_6t_3 inst_cell_127_69 ( BL69, BLN69, WL127);
sram_cell_6t_3 inst_cell_127_68 ( BL68, BLN68, WL127);
sram_cell_6t_3 inst_cell_127_67 ( BL67, BLN67, WL127);
sram_cell_6t_3 inst_cell_127_66 ( BL66, BLN66, WL127);
sram_cell_6t_3 inst_cell_127_65 ( BL65, BLN65, WL127);
sram_cell_6t_3 inst_cell_127_64 ( BL64, BLN64, WL127);
sram_cell_6t_3 inst_cell_127_109 ( BL109, BLN109, WL127);
sram_cell_6t_3 inst_cell_127_108 ( BL108, BLN108, WL127);
sram_cell_6t_3 inst_cell_127_107 ( BL107, BLN107, WL127);
sram_cell_6t_3 inst_cell_127_106 ( BL106, BLN106, WL127);
sram_cell_6t_3 inst_cell_127_105 ( BL105, BLN105, WL127);
sram_cell_6t_3 inst_cell_127_104 ( BL104, BLN104, WL127);
sram_cell_6t_3 inst_cell_127_103 ( BL103, BLN103, WL127);
sram_cell_6t_3 inst_cell_127_102 ( BL102, BLN102, WL127);
sram_cell_6t_3 inst_cell_127_101 ( BL101, BLN101, WL127);
sram_cell_6t_3 inst_cell_127_100 ( BL100, BLN100, WL127);
sram_cell_6t_3 inst_cell_127_99 ( BL99, BLN99, WL127);
sram_cell_6t_3 inst_cell_127_98 ( BL98, BLN98, WL127);
sram_cell_6t_3 inst_cell_127_97 ( BL97, BLN97, WL127);
sram_cell_6t_3 inst_cell_127_96 ( BL96, BLN96, WL127);
sram_cell_6t_3 inst_cell_127_95 ( BL95, BLN95, WL127);
sram_cell_6t_3 inst_cell_127_94 ( BL94, BLN94, WL127);
sram_cell_6t_3 inst_cell_127_93 ( BL93, BLN93, WL127);
sram_cell_6t_3 inst_cell_127_92 ( BL92, BLN92, WL127);
sram_cell_6t_3 inst_cell_127_91 ( BL91, BLN91, WL127);
sram_cell_6t_3 inst_cell_127_90 ( BL90, BLN90, WL127);
sram_cell_6t_3 inst_cell_127_89 ( BL89, BLN89, WL127);
sram_cell_6t_3 inst_cell_127_88 ( BL88, BLN88, WL127);
sram_cell_6t_3 inst_cell_127_87 ( BL87, BLN87, WL127);
sram_cell_6t_3 inst_cell_127_86 ( BL86, BLN86, WL127);
sram_cell_6t_3 inst_cell_127_85 ( BL85, BLN85, WL127);
sram_cell_6t_3 inst_cell_127_84 ( BL84, BLN84, WL127);
sram_cell_6t_3 inst_cell_127_83 ( BL83, BLN83, WL127);
sram_cell_6t_3 inst_cell_127_82 ( BL82, BLN82, WL127);
sram_cell_6t_3 inst_cell_127_81 ( BL81, BLN81, WL127);
sram_cell_6t_3 inst_cell_127_80 ( BL80, BLN80, WL127);
sram_cell_6t_3 inst_cell_127_63 ( BL63, BLN63, WL127);
sram_cell_6t_3 inst_cell_127_62 ( BL62, BLN62, WL127);
sram_cell_6t_3 inst_cell_127_61 ( BL61, BLN61, WL127);
sram_cell_6t_3 inst_cell_127_60 ( BL60, BLN60, WL127);
sram_cell_6t_3 inst_cell_127_59 ( BL59, BLN59, WL127);
sram_cell_6t_3 inst_cell_127_58 ( BL58, BLN58, WL127);
sram_cell_6t_3 inst_cell_127_57 ( BL57, BLN57, WL127);
sram_cell_6t_3 inst_cell_127_56 ( BL56, BLN56, WL127);
sram_cell_6t_3 inst_cell_127_55 ( BL55, BLN55, WL127);
sram_cell_6t_3 inst_cell_127_54 ( BL54, BLN54, WL127);
sram_cell_6t_3 inst_cell_127_53 ( BL53, BLN53, WL127);
sram_cell_6t_3 inst_cell_127_52 ( BL52, BLN52, WL127);
sram_cell_6t_3 inst_cell_127_51 ( BL51, BLN51, WL127);
sram_cell_6t_3 inst_cell_127_50 ( BL50, BLN50, WL127);
sram_cell_6t_3 inst_cell_127_49 ( BL49, BLN49, WL127);
sram_cell_6t_3 inst_cell_127_48 ( BL48, BLN48, WL127);
sram_cell_6t_3 inst_cell_127_47 ( BL47, BLN47, WL127);
sram_cell_6t_3 inst_cell_127_46 ( BL46, BLN46, WL127);
sram_cell_6t_3 inst_cell_127_45 ( BL45, BLN45, WL127);
sram_cell_6t_3 inst_cell_127_44 ( BL44, BLN44, WL127);
sram_cell_6t_3 inst_cell_127_43 ( BL43, BLN43, WL127);
sram_cell_6t_3 inst_cell_127_42 ( BL42, BLN42, WL127);
sram_cell_6t_3 inst_cell_127_41 ( BL41, BLN41, WL127);
sram_cell_6t_3 inst_cell_127_40 ( BL40, BLN40, WL127);
sram_cell_6t_3 inst_cell_127_39 ( BL39, BLN39, WL127);
sram_cell_6t_3 inst_cell_127_38 ( BL38, BLN38, WL127);
sram_cell_6t_3 inst_cell_127_37 ( BL37, BLN37, WL127);
sram_cell_6t_3 inst_cell_127_36 ( BL36, BLN36, WL127);
sram_cell_6t_3 inst_cell_127_35 ( BL35, BLN35, WL127);
sram_cell_6t_3 inst_cell_127_34 ( BL34, BLN34, WL127);
sram_cell_6t_3 inst_cell_127_33 ( BL33, BLN33, WL127);
sram_cell_6t_3 inst_cell_127_32 ( BL32, BLN32, WL127);
sram_cell_6t_3 inst_cell_127_31 ( BL31, BLN31, WL127);
sram_cell_6t_3 inst_cell_127_30 ( BL30, BLN30, WL127);
sram_cell_6t_3 inst_cell_127_29 ( BL29, BLN29, WL127);
sram_cell_6t_3 inst_cell_127_28 ( BL28, BLN28, WL127);
sram_cell_6t_3 inst_cell_127_27 ( BL27, BLN27, WL127);
sram_cell_6t_3 inst_cell_127_26 ( BL26, BLN26, WL127);
sram_cell_6t_3 inst_cell_127_25 ( BL25, BLN25, WL127);
sram_cell_6t_3 inst_cell_127_24 ( BL24, BLN24, WL127);
sram_cell_6t_3 inst_cell_127_23 ( BL23, BLN23, WL127);
sram_cell_6t_3 inst_cell_127_22 ( BL22, BLN22, WL127);
sram_cell_6t_3 inst_cell_127_21 ( BL21, BLN21, WL127);
sram_cell_6t_3 inst_cell_127_20 ( BL20, BLN20, WL127);
sram_cell_6t_3 inst_cell_127_19 ( BL19, BLN19, WL127);
sram_cell_6t_3 inst_cell_127_18 ( BL18, BLN18, WL127);
sram_cell_6t_3 inst_cell_127_17 ( BL17, BLN17, WL127);
sram_cell_6t_3 inst_cell_127_16 ( BL16, BLN16, WL127);
sram_cell_6t_3 inst_cell_127_15 ( BL15, BLN15, WL127);
sram_cell_6t_3 inst_cell_127_14 ( BL14, BLN14, WL127);
sram_cell_6t_3 inst_cell_127_13 ( BL13, BLN13, WL127);
sram_cell_6t_3 inst_cell_127_12 ( BL12, BLN12, WL127);
sram_cell_6t_3 inst_cell_127_11 ( BL11, BLN11, WL127);
sram_cell_6t_3 inst_cell_127_10 ( BL10, BLN10, WL127);
sram_cell_6t_3 inst_cell_127_9 ( BL9, BLN9, WL127);
sram_cell_6t_3 inst_cell_127_8 ( BL8, BLN8, WL127);
sram_cell_6t_3 inst_cell_127_7 ( BL7, BLN7, WL127);
sram_cell_6t_3 inst_cell_127_6 ( BL6, BLN6, WL127);
sram_cell_6t_3 inst_cell_127_5 ( BL5, BLN5, WL127);
sram_cell_6t_3 inst_cell_127_4 ( BL4, BLN4, WL127);
sram_cell_6t_3 inst_cell_126_127 ( BL127, BLN127, WL126);
sram_cell_6t_3 inst_cell_126_126 ( BL126, BLN126, WL126);
sram_cell_6t_3 inst_cell_126_125 ( BL125, BLN125, WL126);
sram_cell_6t_3 inst_cell_126_124 ( BL124, BLN124, WL126);
sram_cell_6t_3 inst_cell_126_123 ( BL123, BLN123, WL126);
sram_cell_6t_3 inst_cell_126_122 ( BL122, BLN122, WL126);
sram_cell_6t_3 inst_cell_126_121 ( BL121, BLN121, WL126);
sram_cell_6t_3 inst_cell_126_120 ( BL120, BLN120, WL126);
sram_cell_6t_3 inst_cell_126_119 ( BL119, BLN119, WL126);
sram_cell_6t_3 inst_cell_126_118 ( BL118, BLN118, WL126);
sram_cell_6t_3 inst_cell_126_117 ( BL117, BLN117, WL126);
sram_cell_6t_3 inst_cell_126_116 ( BL116, BLN116, WL126);
sram_cell_6t_3 inst_cell_126_115 ( BL115, BLN115, WL126);
sram_cell_6t_3 inst_cell_126_114 ( BL114, BLN114, WL126);
sram_cell_6t_3 inst_cell_126_113 ( BL113, BLN113, WL126);
sram_cell_6t_3 inst_cell_126_112 ( BL112, BLN112, WL126);
sram_cell_6t_3 inst_cell_126_111 ( BL111, BLN111, WL126);
sram_cell_6t_3 inst_cell_126_110 ( BL110, BLN110, WL126);
sram_cell_6t_3 inst_cell_126_109 ( BL109, BLN109, WL126);
sram_cell_6t_3 inst_cell_126_108 ( BL108, BLN108, WL126);
sram_cell_6t_3 inst_cell_126_107 ( BL107, BLN107, WL126);
sram_cell_6t_3 inst_cell_126_106 ( BL106, BLN106, WL126);
sram_cell_6t_3 inst_cell_126_105 ( BL105, BLN105, WL126);
sram_cell_6t_3 inst_cell_126_104 ( BL104, BLN104, WL126);
sram_cell_6t_3 inst_cell_126_103 ( BL103, BLN103, WL126);
sram_cell_6t_3 inst_cell_126_102 ( BL102, BLN102, WL126);
sram_cell_6t_3 inst_cell_126_101 ( BL101, BLN101, WL126);
sram_cell_6t_3 inst_cell_126_100 ( BL100, BLN100, WL126);
sram_cell_6t_3 inst_cell_126_99 ( BL99, BLN99, WL126);
sram_cell_6t_3 inst_cell_126_98 ( BL98, BLN98, WL126);
sram_cell_6t_3 inst_cell_126_97 ( BL97, BLN97, WL126);
sram_cell_6t_3 inst_cell_126_96 ( BL96, BLN96, WL126);
sram_cell_6t_3 inst_cell_126_95 ( BL95, BLN95, WL126);
sram_cell_6t_3 inst_cell_126_94 ( BL94, BLN94, WL126);
sram_cell_6t_3 inst_cell_126_93 ( BL93, BLN93, WL126);
sram_cell_6t_3 inst_cell_126_92 ( BL92, BLN92, WL126);
sram_cell_6t_3 inst_cell_126_91 ( BL91, BLN91, WL126);
sram_cell_6t_3 inst_cell_126_90 ( BL90, BLN90, WL126);
sram_cell_6t_3 inst_cell_126_89 ( BL89, BLN89, WL126);
sram_cell_6t_3 inst_cell_126_88 ( BL88, BLN88, WL126);
sram_cell_6t_3 inst_cell_126_87 ( BL87, BLN87, WL126);
sram_cell_6t_3 inst_cell_126_86 ( BL86, BLN86, WL126);
sram_cell_6t_3 inst_cell_126_85 ( BL85, BLN85, WL126);
sram_cell_6t_3 inst_cell_126_84 ( BL84, BLN84, WL126);
sram_cell_6t_3 inst_cell_126_83 ( BL83, BLN83, WL126);
sram_cell_6t_3 inst_cell_126_82 ( BL82, BLN82, WL126);
sram_cell_6t_3 inst_cell_126_81 ( BL81, BLN81, WL126);
sram_cell_6t_3 inst_cell_126_80 ( BL80, BLN80, WL126);
sram_cell_6t_3 inst_cell_126_79 ( BL79, BLN79, WL126);
sram_cell_6t_3 inst_cell_126_78 ( BL78, BLN78, WL126);
sram_cell_6t_3 inst_cell_126_77 ( BL77, BLN77, WL126);
sram_cell_6t_3 inst_cell_126_76 ( BL76, BLN76, WL126);
sram_cell_6t_3 inst_cell_126_75 ( BL75, BLN75, WL126);
sram_cell_6t_3 inst_cell_126_74 ( BL74, BLN74, WL126);
sram_cell_6t_3 inst_cell_126_73 ( BL73, BLN73, WL126);
sram_cell_6t_3 inst_cell_126_72 ( BL72, BLN72, WL126);
sram_cell_6t_3 inst_cell_126_71 ( BL71, BLN71, WL126);
sram_cell_6t_3 inst_cell_126_70 ( BL70, BLN70, WL126);
sram_cell_6t_3 inst_cell_126_69 ( BL69, BLN69, WL126);
sram_cell_6t_3 inst_cell_126_68 ( BL68, BLN68, WL126);
sram_cell_6t_3 inst_cell_126_67 ( BL67, BLN67, WL126);
sram_cell_6t_3 inst_cell_126_66 ( BL66, BLN66, WL126);
sram_cell_6t_3 inst_cell_126_65 ( BL65, BLN65, WL126);
sram_cell_6t_3 inst_cell_126_64 ( BL64, BLN64, WL126);
sram_cell_6t_3 inst_cell_126_63 ( BL63, BLN63, WL126);
sram_cell_6t_3 inst_cell_126_62 ( BL62, BLN62, WL126);
sram_cell_6t_3 inst_cell_126_61 ( BL61, BLN61, WL126);
sram_cell_6t_3 inst_cell_126_60 ( BL60, BLN60, WL126);
sram_cell_6t_3 inst_cell_126_59 ( BL59, BLN59, WL126);
sram_cell_6t_3 inst_cell_126_58 ( BL58, BLN58, WL126);
sram_cell_6t_3 inst_cell_126_57 ( BL57, BLN57, WL126);
sram_cell_6t_3 inst_cell_126_56 ( BL56, BLN56, WL126);
sram_cell_6t_3 inst_cell_126_55 ( BL55, BLN55, WL126);
sram_cell_6t_3 inst_cell_126_54 ( BL54, BLN54, WL126);
sram_cell_6t_3 inst_cell_126_53 ( BL53, BLN53, WL126);
sram_cell_6t_3 inst_cell_126_52 ( BL52, BLN52, WL126);
sram_cell_6t_3 inst_cell_126_51 ( BL51, BLN51, WL126);
sram_cell_6t_3 inst_cell_126_50 ( BL50, BLN50, WL126);
sram_cell_6t_3 inst_cell_126_49 ( BL49, BLN49, WL126);
sram_cell_6t_3 inst_cell_126_48 ( BL48, BLN48, WL126);
sram_cell_6t_3 inst_cell_126_47 ( BL47, BLN47, WL126);
sram_cell_6t_3 inst_cell_126_46 ( BL46, BLN46, WL126);
sram_cell_6t_3 inst_cell_126_45 ( BL45, BLN45, WL126);
sram_cell_6t_3 inst_cell_126_44 ( BL44, BLN44, WL126);
sram_cell_6t_3 inst_cell_126_43 ( BL43, BLN43, WL126);
sram_cell_6t_3 inst_cell_126_42 ( BL42, BLN42, WL126);
sram_cell_6t_3 inst_cell_126_41 ( BL41, BLN41, WL126);
sram_cell_6t_3 inst_cell_126_40 ( BL40, BLN40, WL126);
sram_cell_6t_3 inst_cell_126_15 ( BL15, BLN15, WL126);
sram_cell_6t_3 inst_cell_126_14 ( BL14, BLN14, WL126);
sram_cell_6t_3 inst_cell_126_13 ( BL13, BLN13, WL126);
sram_cell_6t_3 inst_cell_126_12 ( BL12, BLN12, WL126);
sram_cell_6t_3 inst_cell_126_11 ( BL11, BLN11, WL126);
sram_cell_6t_3 inst_cell_126_10 ( BL10, BLN10, WL126);
sram_cell_6t_3 inst_cell_126_9 ( BL9, BLN9, WL126);
sram_cell_6t_3 inst_cell_126_8 ( BL8, BLN8, WL126);
sram_cell_6t_3 inst_cell_126_7 ( BL7, BLN7, WL126);
sram_cell_6t_3 inst_cell_126_6 ( BL6, BLN6, WL126);
sram_cell_6t_3 inst_cell_126_5 ( BL5, BLN5, WL126);
sram_cell_6t_3 inst_cell_126_4 ( BL4, BLN4, WL126);
sram_cell_6t_3 inst_cell_126_3 ( BL3, BLN3, WL126);
sram_cell_6t_3 inst_cell_126_2 ( BL2, BLN2, WL126);
sram_cell_6t_3 inst_cell_126_1 ( BL1, BLN1, WL126);
sram_cell_6t_3 inst_cell_126_0 ( BL0, BLN0, WL126);
sram_cell_6t_3 inst_cell_126_39 ( BL39, BLN39, WL126);
sram_cell_6t_3 inst_cell_126_38 ( BL38, BLN38, WL126);
sram_cell_6t_3 inst_cell_126_37 ( BL37, BLN37, WL126);
sram_cell_6t_3 inst_cell_126_36 ( BL36, BLN36, WL126);
sram_cell_6t_3 inst_cell_126_35 ( BL35, BLN35, WL126);
sram_cell_6t_3 inst_cell_126_34 ( BL34, BLN34, WL126);
sram_cell_6t_3 inst_cell_126_33 ( BL33, BLN33, WL126);
sram_cell_6t_3 inst_cell_126_32 ( BL32, BLN32, WL126);
sram_cell_6t_3 inst_cell_126_31 ( BL31, BLN31, WL126);
sram_cell_6t_3 inst_cell_126_30 ( BL30, BLN30, WL126);
sram_cell_6t_3 inst_cell_126_29 ( BL29, BLN29, WL126);
sram_cell_6t_3 inst_cell_126_28 ( BL28, BLN28, WL126);
sram_cell_6t_3 inst_cell_126_27 ( BL27, BLN27, WL126);
sram_cell_6t_3 inst_cell_126_26 ( BL26, BLN26, WL126);
sram_cell_6t_3 inst_cell_126_25 ( BL25, BLN25, WL126);
sram_cell_6t_3 inst_cell_126_24 ( BL24, BLN24, WL126);
sram_cell_6t_3 inst_cell_126_23 ( BL23, BLN23, WL126);
sram_cell_6t_3 inst_cell_126_22 ( BL22, BLN22, WL126);
sram_cell_6t_3 inst_cell_126_21 ( BL21, BLN21, WL126);
sram_cell_6t_3 inst_cell_126_20 ( BL20, BLN20, WL126);
sram_cell_6t_3 inst_cell_126_19 ( BL19, BLN19, WL126);
sram_cell_6t_3 inst_cell_126_18 ( BL18, BLN18, WL126);
sram_cell_6t_3 inst_cell_126_17 ( BL17, BLN17, WL126);
sram_cell_6t_3 inst_cell_126_16 ( BL16, BLN16, WL126);
sram_cell_6t_3 inst_cell_125_127 ( BL127, BLN127, WL125);
sram_cell_6t_3 inst_cell_125_126 ( BL126, BLN126, WL125);
sram_cell_6t_3 inst_cell_125_125 ( BL125, BLN125, WL125);
sram_cell_6t_3 inst_cell_125_124 ( BL124, BLN124, WL125);
sram_cell_6t_3 inst_cell_125_123 ( BL123, BLN123, WL125);
sram_cell_6t_3 inst_cell_125_122 ( BL122, BLN122, WL125);
sram_cell_6t_3 inst_cell_125_121 ( BL121, BLN121, WL125);
sram_cell_6t_3 inst_cell_125_120 ( BL120, BLN120, WL125);
sram_cell_6t_3 inst_cell_125_119 ( BL119, BLN119, WL125);
sram_cell_6t_3 inst_cell_125_118 ( BL118, BLN118, WL125);
sram_cell_6t_3 inst_cell_125_117 ( BL117, BLN117, WL125);
sram_cell_6t_3 inst_cell_125_116 ( BL116, BLN116, WL125);
sram_cell_6t_3 inst_cell_125_115 ( BL115, BLN115, WL125);
sram_cell_6t_3 inst_cell_125_114 ( BL114, BLN114, WL125);
sram_cell_6t_3 inst_cell_125_113 ( BL113, BLN113, WL125);
sram_cell_6t_3 inst_cell_125_112 ( BL112, BLN112, WL125);
sram_cell_6t_3 inst_cell_125_111 ( BL111, BLN111, WL125);
sram_cell_6t_3 inst_cell_125_110 ( BL110, BLN110, WL125);
sram_cell_6t_3 inst_cell_125_109 ( BL109, BLN109, WL125);
sram_cell_6t_3 inst_cell_125_108 ( BL108, BLN108, WL125);
sram_cell_6t_3 inst_cell_125_107 ( BL107, BLN107, WL125);
sram_cell_6t_3 inst_cell_125_106 ( BL106, BLN106, WL125);
sram_cell_6t_3 inst_cell_125_105 ( BL105, BLN105, WL125);
sram_cell_6t_3 inst_cell_125_104 ( BL104, BLN104, WL125);
sram_cell_6t_3 inst_cell_125_103 ( BL103, BLN103, WL125);
sram_cell_6t_3 inst_cell_125_102 ( BL102, BLN102, WL125);
sram_cell_6t_3 inst_cell_125_101 ( BL101, BLN101, WL125);
sram_cell_6t_3 inst_cell_125_100 ( BL100, BLN100, WL125);
sram_cell_6t_3 inst_cell_125_99 ( BL99, BLN99, WL125);
sram_cell_6t_3 inst_cell_125_98 ( BL98, BLN98, WL125);
sram_cell_6t_3 inst_cell_125_97 ( BL97, BLN97, WL125);
sram_cell_6t_3 inst_cell_125_96 ( BL96, BLN96, WL125);
sram_cell_6t_3 inst_cell_125_95 ( BL95, BLN95, WL125);
sram_cell_6t_3 inst_cell_125_94 ( BL94, BLN94, WL125);
sram_cell_6t_3 inst_cell_125_93 ( BL93, BLN93, WL125);
sram_cell_6t_3 inst_cell_125_92 ( BL92, BLN92, WL125);
sram_cell_6t_3 inst_cell_125_91 ( BL91, BLN91, WL125);
sram_cell_6t_3 inst_cell_125_90 ( BL90, BLN90, WL125);
sram_cell_6t_3 inst_cell_125_89 ( BL89, BLN89, WL125);
sram_cell_6t_3 inst_cell_125_88 ( BL88, BLN88, WL125);
sram_cell_6t_3 inst_cell_125_87 ( BL87, BLN87, WL125);
sram_cell_6t_3 inst_cell_125_86 ( BL86, BLN86, WL125);
sram_cell_6t_3 inst_cell_125_85 ( BL85, BLN85, WL125);
sram_cell_6t_3 inst_cell_125_84 ( BL84, BLN84, WL125);
sram_cell_6t_3 inst_cell_125_83 ( BL83, BLN83, WL125);
sram_cell_6t_3 inst_cell_125_82 ( BL82, BLN82, WL125);
sram_cell_6t_3 inst_cell_125_81 ( BL81, BLN81, WL125);
sram_cell_6t_3 inst_cell_125_80 ( BL80, BLN80, WL125);
sram_cell_6t_3 inst_cell_125_79 ( BL79, BLN79, WL125);
sram_cell_6t_3 inst_cell_125_78 ( BL78, BLN78, WL125);
sram_cell_6t_3 inst_cell_125_77 ( BL77, BLN77, WL125);
sram_cell_6t_3 inst_cell_125_76 ( BL76, BLN76, WL125);
sram_cell_6t_3 inst_cell_125_75 ( BL75, BLN75, WL125);
sram_cell_6t_3 inst_cell_125_74 ( BL74, BLN74, WL125);
sram_cell_6t_3 inst_cell_125_73 ( BL73, BLN73, WL125);
sram_cell_6t_3 inst_cell_125_72 ( BL72, BLN72, WL125);
sram_cell_6t_3 inst_cell_125_71 ( BL71, BLN71, WL125);
sram_cell_6t_3 inst_cell_125_70 ( BL70, BLN70, WL125);
sram_cell_6t_3 inst_cell_125_69 ( BL69, BLN69, WL125);
sram_cell_6t_3 inst_cell_125_68 ( BL68, BLN68, WL125);
sram_cell_6t_3 inst_cell_125_67 ( BL67, BLN67, WL125);
sram_cell_6t_3 inst_cell_125_66 ( BL66, BLN66, WL125);
sram_cell_6t_3 inst_cell_125_65 ( BL65, BLN65, WL125);
sram_cell_6t_3 inst_cell_125_64 ( BL64, BLN64, WL125);
sram_cell_6t_3 inst_cell_125_63 ( BL63, BLN63, WL125);
sram_cell_6t_3 inst_cell_125_62 ( BL62, BLN62, WL125);
sram_cell_6t_3 inst_cell_125_61 ( BL61, BLN61, WL125);
sram_cell_6t_3 inst_cell_125_60 ( BL60, BLN60, WL125);
sram_cell_6t_3 inst_cell_125_59 ( BL59, BLN59, WL125);
sram_cell_6t_3 inst_cell_125_58 ( BL58, BLN58, WL125);
sram_cell_6t_3 inst_cell_125_57 ( BL57, BLN57, WL125);
sram_cell_6t_3 inst_cell_125_56 ( BL56, BLN56, WL125);
sram_cell_6t_3 inst_cell_125_55 ( BL55, BLN55, WL125);
sram_cell_6t_3 inst_cell_125_54 ( BL54, BLN54, WL125);
sram_cell_6t_3 inst_cell_125_53 ( BL53, BLN53, WL125);
sram_cell_6t_3 inst_cell_125_52 ( BL52, BLN52, WL125);
sram_cell_6t_3 inst_cell_125_51 ( BL51, BLN51, WL125);
sram_cell_6t_3 inst_cell_125_50 ( BL50, BLN50, WL125);
sram_cell_6t_3 inst_cell_125_49 ( BL49, BLN49, WL125);
sram_cell_6t_3 inst_cell_125_48 ( BL48, BLN48, WL125);
sram_cell_6t_3 inst_cell_125_47 ( BL47, BLN47, WL125);
sram_cell_6t_3 inst_cell_125_46 ( BL46, BLN46, WL125);
sram_cell_6t_3 inst_cell_125_45 ( BL45, BLN45, WL125);
sram_cell_6t_3 inst_cell_125_44 ( BL44, BLN44, WL125);
sram_cell_6t_3 inst_cell_125_43 ( BL43, BLN43, WL125);
sram_cell_6t_3 inst_cell_125_42 ( BL42, BLN42, WL125);
sram_cell_6t_3 inst_cell_125_41 ( BL41, BLN41, WL125);
sram_cell_6t_3 inst_cell_125_40 ( BL40, BLN40, WL125);
sram_cell_6t_3 inst_cell_125_39 ( BL39, BLN39, WL125);
sram_cell_6t_3 inst_cell_125_38 ( BL38, BLN38, WL125);
sram_cell_6t_3 inst_cell_125_37 ( BL37, BLN37, WL125);
sram_cell_6t_3 inst_cell_125_36 ( BL36, BLN36, WL125);
sram_cell_6t_3 inst_cell_125_35 ( BL35, BLN35, WL125);
sram_cell_6t_3 inst_cell_125_34 ( BL34, BLN34, WL125);
sram_cell_6t_3 inst_cell_125_33 ( BL33, BLN33, WL125);
sram_cell_6t_3 inst_cell_125_32 ( BL32, BLN32, WL125);
sram_cell_6t_3 inst_cell_125_31 ( BL31, BLN31, WL125);
sram_cell_6t_3 inst_cell_125_30 ( BL30, BLN30, WL125);
sram_cell_6t_3 inst_cell_125_29 ( BL29, BLN29, WL125);
sram_cell_6t_3 inst_cell_125_28 ( BL28, BLN28, WL125);
sram_cell_6t_3 inst_cell_125_27 ( BL27, BLN27, WL125);
sram_cell_6t_3 inst_cell_125_26 ( BL26, BLN26, WL125);
sram_cell_6t_3 inst_cell_125_25 ( BL25, BLN25, WL125);
sram_cell_6t_3 inst_cell_125_24 ( BL24, BLN24, WL125);
sram_cell_6t_3 inst_cell_125_23 ( BL23, BLN23, WL125);
sram_cell_6t_3 inst_cell_125_22 ( BL22, BLN22, WL125);
sram_cell_6t_3 inst_cell_125_21 ( BL21, BLN21, WL125);
sram_cell_6t_3 inst_cell_125_20 ( BL20, BLN20, WL125);
sram_cell_6t_3 inst_cell_125_19 ( BL19, BLN19, WL125);
sram_cell_6t_3 inst_cell_125_18 ( BL18, BLN18, WL125);
sram_cell_6t_3 inst_cell_125_17 ( BL17, BLN17, WL125);
sram_cell_6t_3 inst_cell_125_16 ( BL16, BLN16, WL125);
sram_cell_6t_3 inst_cell_125_15 ( BL15, BLN15, WL125);
sram_cell_6t_3 inst_cell_125_14 ( BL14, BLN14, WL125);
sram_cell_6t_3 inst_cell_125_13 ( BL13, BLN13, WL125);
sram_cell_6t_3 inst_cell_125_12 ( BL12, BLN12, WL125);
sram_cell_6t_3 inst_cell_125_11 ( BL11, BLN11, WL125);
sram_cell_6t_3 inst_cell_125_10 ( BL10, BLN10, WL125);
sram_cell_6t_3 inst_cell_125_9 ( BL9, BLN9, WL125);
sram_cell_6t_3 inst_cell_125_8 ( BL8, BLN8, WL125);
sram_cell_6t_3 inst_cell_125_7 ( BL7, BLN7, WL125);
sram_cell_6t_3 inst_cell_125_6 ( BL6, BLN6, WL125);
sram_cell_6t_3 inst_cell_125_5 ( BL5, BLN5, WL125);
sram_cell_6t_3 inst_cell_125_4 ( BL4, BLN4, WL125);
sram_cell_6t_3 inst_cell_125_3 ( BL3, BLN3, WL125);
sram_cell_6t_3 inst_cell_125_2 ( BL2, BLN2, WL125);
sram_cell_6t_3 inst_cell_125_1 ( BL1, BLN1, WL125);
sram_cell_6t_3 inst_cell_125_0 ( BL0, BLN0, WL125);
sram_cell_6t_3 inst_cell_124_127 ( BL127, BLN127, WL124);
sram_cell_6t_3 inst_cell_124_126 ( BL126, BLN126, WL124);
sram_cell_6t_3 inst_cell_124_125 ( BL125, BLN125, WL124);
sram_cell_6t_3 inst_cell_124_124 ( BL124, BLN124, WL124);
sram_cell_6t_3 inst_cell_124_123 ( BL123, BLN123, WL124);
sram_cell_6t_3 inst_cell_124_122 ( BL122, BLN122, WL124);
sram_cell_6t_3 inst_cell_124_121 ( BL121, BLN121, WL124);
sram_cell_6t_3 inst_cell_124_120 ( BL120, BLN120, WL124);
sram_cell_6t_3 inst_cell_124_119 ( BL119, BLN119, WL124);
sram_cell_6t_3 inst_cell_124_118 ( BL118, BLN118, WL124);
sram_cell_6t_3 inst_cell_124_117 ( BL117, BLN117, WL124);
sram_cell_6t_3 inst_cell_124_116 ( BL116, BLN116, WL124);
sram_cell_6t_3 inst_cell_124_115 ( BL115, BLN115, WL124);
sram_cell_6t_3 inst_cell_124_114 ( BL114, BLN114, WL124);
sram_cell_6t_3 inst_cell_124_113 ( BL113, BLN113, WL124);
sram_cell_6t_3 inst_cell_124_112 ( BL112, BLN112, WL124);
sram_cell_6t_3 inst_cell_124_111 ( BL111, BLN111, WL124);
sram_cell_6t_3 inst_cell_124_110 ( BL110, BLN110, WL124);
sram_cell_6t_3 inst_cell_124_109 ( BL109, BLN109, WL124);
sram_cell_6t_3 inst_cell_124_108 ( BL108, BLN108, WL124);
sram_cell_6t_3 inst_cell_124_107 ( BL107, BLN107, WL124);
sram_cell_6t_3 inst_cell_124_106 ( BL106, BLN106, WL124);
sram_cell_6t_3 inst_cell_124_105 ( BL105, BLN105, WL124);
sram_cell_6t_3 inst_cell_124_104 ( BL104, BLN104, WL124);
sram_cell_6t_3 inst_cell_124_103 ( BL103, BLN103, WL124);
sram_cell_6t_3 inst_cell_124_102 ( BL102, BLN102, WL124);
sram_cell_6t_3 inst_cell_124_101 ( BL101, BLN101, WL124);
sram_cell_6t_3 inst_cell_124_100 ( BL100, BLN100, WL124);
sram_cell_6t_3 inst_cell_124_99 ( BL99, BLN99, WL124);
sram_cell_6t_3 inst_cell_124_98 ( BL98, BLN98, WL124);
sram_cell_6t_3 inst_cell_124_97 ( BL97, BLN97, WL124);
sram_cell_6t_3 inst_cell_124_96 ( BL96, BLN96, WL124);
sram_cell_6t_3 inst_cell_124_95 ( BL95, BLN95, WL124);
sram_cell_6t_3 inst_cell_124_94 ( BL94, BLN94, WL124);
sram_cell_6t_3 inst_cell_124_93 ( BL93, BLN93, WL124);
sram_cell_6t_3 inst_cell_124_92 ( BL92, BLN92, WL124);
sram_cell_6t_3 inst_cell_124_91 ( BL91, BLN91, WL124);
sram_cell_6t_3 inst_cell_124_90 ( BL90, BLN90, WL124);
sram_cell_6t_3 inst_cell_124_89 ( BL89, BLN89, WL124);
sram_cell_6t_3 inst_cell_124_88 ( BL88, BLN88, WL124);
sram_cell_6t_3 inst_cell_124_87 ( BL87, BLN87, WL124);
sram_cell_6t_3 inst_cell_124_86 ( BL86, BLN86, WL124);
sram_cell_6t_3 inst_cell_124_85 ( BL85, BLN85, WL124);
sram_cell_6t_3 inst_cell_124_84 ( BL84, BLN84, WL124);
sram_cell_6t_3 inst_cell_124_83 ( BL83, BLN83, WL124);
sram_cell_6t_3 inst_cell_124_82 ( BL82, BLN82, WL124);
sram_cell_6t_3 inst_cell_124_81 ( BL81, BLN81, WL124);
sram_cell_6t_3 inst_cell_124_80 ( BL80, BLN80, WL124);
sram_cell_6t_3 inst_cell_124_79 ( BL79, BLN79, WL124);
sram_cell_6t_3 inst_cell_124_78 ( BL78, BLN78, WL124);
sram_cell_6t_3 inst_cell_124_77 ( BL77, BLN77, WL124);
sram_cell_6t_3 inst_cell_124_76 ( BL76, BLN76, WL124);
sram_cell_6t_3 inst_cell_124_75 ( BL75, BLN75, WL124);
sram_cell_6t_3 inst_cell_124_74 ( BL74, BLN74, WL124);
sram_cell_6t_3 inst_cell_124_73 ( BL73, BLN73, WL124);
sram_cell_6t_3 inst_cell_124_72 ( BL72, BLN72, WL124);
sram_cell_6t_3 inst_cell_124_71 ( BL71, BLN71, WL124);
sram_cell_6t_3 inst_cell_124_70 ( BL70, BLN70, WL124);
sram_cell_6t_3 inst_cell_124_69 ( BL69, BLN69, WL124);
sram_cell_6t_3 inst_cell_124_68 ( BL68, BLN68, WL124);
sram_cell_6t_3 inst_cell_124_67 ( BL67, BLN67, WL124);
sram_cell_6t_3 inst_cell_124_66 ( BL66, BLN66, WL124);
sram_cell_6t_3 inst_cell_124_65 ( BL65, BLN65, WL124);
sram_cell_6t_3 inst_cell_124_64 ( BL64, BLN64, WL124);
sram_cell_6t_3 inst_cell_124_63 ( BL63, BLN63, WL124);
sram_cell_6t_3 inst_cell_124_62 ( BL62, BLN62, WL124);
sram_cell_6t_3 inst_cell_124_61 ( BL61, BLN61, WL124);
sram_cell_6t_3 inst_cell_124_60 ( BL60, BLN60, WL124);
sram_cell_6t_3 inst_cell_124_59 ( BL59, BLN59, WL124);
sram_cell_6t_3 inst_cell_124_58 ( BL58, BLN58, WL124);
sram_cell_6t_3 inst_cell_124_57 ( BL57, BLN57, WL124);
sram_cell_6t_3 inst_cell_124_56 ( BL56, BLN56, WL124);
sram_cell_6t_3 inst_cell_124_55 ( BL55, BLN55, WL124);
sram_cell_6t_3 inst_cell_124_54 ( BL54, BLN54, WL124);
sram_cell_6t_3 inst_cell_124_53 ( BL53, BLN53, WL124);
sram_cell_6t_3 inst_cell_124_52 ( BL52, BLN52, WL124);
sram_cell_6t_3 inst_cell_124_51 ( BL51, BLN51, WL124);
sram_cell_6t_3 inst_cell_124_50 ( BL50, BLN50, WL124);
sram_cell_6t_3 inst_cell_124_49 ( BL49, BLN49, WL124);
sram_cell_6t_3 inst_cell_124_48 ( BL48, BLN48, WL124);
sram_cell_6t_3 inst_cell_124_47 ( BL47, BLN47, WL124);
sram_cell_6t_3 inst_cell_124_46 ( BL46, BLN46, WL124);
sram_cell_6t_3 inst_cell_124_45 ( BL45, BLN45, WL124);
sram_cell_6t_3 inst_cell_124_44 ( BL44, BLN44, WL124);
sram_cell_6t_3 inst_cell_124_43 ( BL43, BLN43, WL124);
sram_cell_6t_3 inst_cell_124_42 ( BL42, BLN42, WL124);
sram_cell_6t_3 inst_cell_124_41 ( BL41, BLN41, WL124);
sram_cell_6t_3 inst_cell_124_40 ( BL40, BLN40, WL124);
sram_cell_6t_3 inst_cell_124_39 ( BL39, BLN39, WL124);
sram_cell_6t_3 inst_cell_124_38 ( BL38, BLN38, WL124);
sram_cell_6t_3 inst_cell_124_37 ( BL37, BLN37, WL124);
sram_cell_6t_3 inst_cell_124_36 ( BL36, BLN36, WL124);
sram_cell_6t_3 inst_cell_124_35 ( BL35, BLN35, WL124);
sram_cell_6t_3 inst_cell_124_34 ( BL34, BLN34, WL124);
sram_cell_6t_3 inst_cell_124_33 ( BL33, BLN33, WL124);
sram_cell_6t_3 inst_cell_124_32 ( BL32, BLN32, WL124);
sram_cell_6t_3 inst_cell_124_31 ( BL31, BLN31, WL124);
sram_cell_6t_3 inst_cell_124_30 ( BL30, BLN30, WL124);
sram_cell_6t_3 inst_cell_124_29 ( BL29, BLN29, WL124);
sram_cell_6t_3 inst_cell_124_28 ( BL28, BLN28, WL124);
sram_cell_6t_3 inst_cell_124_27 ( BL27, BLN27, WL124);
sram_cell_6t_3 inst_cell_124_26 ( BL26, BLN26, WL124);
sram_cell_6t_3 inst_cell_124_25 ( BL25, BLN25, WL124);
sram_cell_6t_3 inst_cell_124_24 ( BL24, BLN24, WL124);
sram_cell_6t_3 inst_cell_124_23 ( BL23, BLN23, WL124);
sram_cell_6t_3 inst_cell_124_22 ( BL22, BLN22, WL124);
sram_cell_6t_3 inst_cell_124_21 ( BL21, BLN21, WL124);
sram_cell_6t_3 inst_cell_124_20 ( BL20, BLN20, WL124);
sram_cell_6t_3 inst_cell_124_19 ( BL19, BLN19, WL124);
sram_cell_6t_3 inst_cell_124_18 ( BL18, BLN18, WL124);
sram_cell_6t_3 inst_cell_124_17 ( BL17, BLN17, WL124);
sram_cell_6t_3 inst_cell_124_16 ( BL16, BLN16, WL124);
sram_cell_6t_3 inst_cell_124_15 ( BL15, BLN15, WL124);
sram_cell_6t_3 inst_cell_124_14 ( BL14, BLN14, WL124);
sram_cell_6t_3 inst_cell_124_13 ( BL13, BLN13, WL124);
sram_cell_6t_3 inst_cell_124_12 ( BL12, BLN12, WL124);
sram_cell_6t_3 inst_cell_124_11 ( BL11, BLN11, WL124);
sram_cell_6t_3 inst_cell_124_10 ( BL10, BLN10, WL124);
sram_cell_6t_3 inst_cell_124_9 ( BL9, BLN9, WL124);
sram_cell_6t_3 inst_cell_124_8 ( BL8, BLN8, WL124);
sram_cell_6t_3 inst_cell_124_7 ( BL7, BLN7, WL124);
sram_cell_6t_3 inst_cell_124_6 ( BL6, BLN6, WL124);
sram_cell_6t_3 inst_cell_124_5 ( BL5, BLN5, WL124);
sram_cell_6t_3 inst_cell_124_4 ( BL4, BLN4, WL124);
sram_cell_6t_3 inst_cell_124_3 ( BL3, BLN3, WL124);
sram_cell_6t_3 inst_cell_124_2 ( BL2, BLN2, WL124);
sram_cell_6t_3 inst_cell_124_1 ( BL1, BLN1, WL124);
sram_cell_6t_3 inst_cell_124_0 ( BL0, BLN0, WL124);
sram_cell_6t_3 inst_cell_123_127 ( BL127, BLN127, WL123);
sram_cell_6t_3 inst_cell_123_126 ( BL126, BLN126, WL123);
sram_cell_6t_3 inst_cell_123_125 ( BL125, BLN125, WL123);
sram_cell_6t_3 inst_cell_123_124 ( BL124, BLN124, WL123);
sram_cell_6t_3 inst_cell_123_123 ( BL123, BLN123, WL123);
sram_cell_6t_3 inst_cell_123_122 ( BL122, BLN122, WL123);
sram_cell_6t_3 inst_cell_123_121 ( BL121, BLN121, WL123);
sram_cell_6t_3 inst_cell_123_120 ( BL120, BLN120, WL123);
sram_cell_6t_3 inst_cell_123_119 ( BL119, BLN119, WL123);
sram_cell_6t_3 inst_cell_123_118 ( BL118, BLN118, WL123);
sram_cell_6t_3 inst_cell_123_117 ( BL117, BLN117, WL123);
sram_cell_6t_3 inst_cell_123_116 ( BL116, BLN116, WL123);
sram_cell_6t_3 inst_cell_123_115 ( BL115, BLN115, WL123);
sram_cell_6t_3 inst_cell_123_114 ( BL114, BLN114, WL123);
sram_cell_6t_3 inst_cell_123_113 ( BL113, BLN113, WL123);
sram_cell_6t_3 inst_cell_123_112 ( BL112, BLN112, WL123);
sram_cell_6t_3 inst_cell_123_111 ( BL111, BLN111, WL123);
sram_cell_6t_3 inst_cell_123_110 ( BL110, BLN110, WL123);
sram_cell_6t_3 inst_cell_123_109 ( BL109, BLN109, WL123);
sram_cell_6t_3 inst_cell_123_108 ( BL108, BLN108, WL123);
sram_cell_6t_3 inst_cell_123_107 ( BL107, BLN107, WL123);
sram_cell_6t_3 inst_cell_123_106 ( BL106, BLN106, WL123);
sram_cell_6t_3 inst_cell_123_105 ( BL105, BLN105, WL123);
sram_cell_6t_3 inst_cell_123_104 ( BL104, BLN104, WL123);
sram_cell_6t_3 inst_cell_123_103 ( BL103, BLN103, WL123);
sram_cell_6t_3 inst_cell_123_102 ( BL102, BLN102, WL123);
sram_cell_6t_3 inst_cell_123_101 ( BL101, BLN101, WL123);
sram_cell_6t_3 inst_cell_123_100 ( BL100, BLN100, WL123);
sram_cell_6t_3 inst_cell_123_99 ( BL99, BLN99, WL123);
sram_cell_6t_3 inst_cell_123_98 ( BL98, BLN98, WL123);
sram_cell_6t_3 inst_cell_123_97 ( BL97, BLN97, WL123);
sram_cell_6t_3 inst_cell_123_96 ( BL96, BLN96, WL123);
sram_cell_6t_3 inst_cell_123_95 ( BL95, BLN95, WL123);
sram_cell_6t_3 inst_cell_123_94 ( BL94, BLN94, WL123);
sram_cell_6t_3 inst_cell_123_93 ( BL93, BLN93, WL123);
sram_cell_6t_3 inst_cell_123_92 ( BL92, BLN92, WL123);
sram_cell_6t_3 inst_cell_123_91 ( BL91, BLN91, WL123);
sram_cell_6t_3 inst_cell_123_90 ( BL90, BLN90, WL123);
sram_cell_6t_3 inst_cell_123_89 ( BL89, BLN89, WL123);
sram_cell_6t_3 inst_cell_123_88 ( BL88, BLN88, WL123);
sram_cell_6t_3 inst_cell_123_87 ( BL87, BLN87, WL123);
sram_cell_6t_3 inst_cell_123_86 ( BL86, BLN86, WL123);
sram_cell_6t_3 inst_cell_123_85 ( BL85, BLN85, WL123);
sram_cell_6t_3 inst_cell_123_84 ( BL84, BLN84, WL123);
sram_cell_6t_3 inst_cell_123_83 ( BL83, BLN83, WL123);
sram_cell_6t_3 inst_cell_123_82 ( BL82, BLN82, WL123);
sram_cell_6t_3 inst_cell_123_81 ( BL81, BLN81, WL123);
sram_cell_6t_3 inst_cell_123_80 ( BL80, BLN80, WL123);
sram_cell_6t_3 inst_cell_123_79 ( BL79, BLN79, WL123);
sram_cell_6t_3 inst_cell_123_78 ( BL78, BLN78, WL123);
sram_cell_6t_3 inst_cell_123_77 ( BL77, BLN77, WL123);
sram_cell_6t_3 inst_cell_123_76 ( BL76, BLN76, WL123);
sram_cell_6t_3 inst_cell_123_75 ( BL75, BLN75, WL123);
sram_cell_6t_3 inst_cell_123_74 ( BL74, BLN74, WL123);
sram_cell_6t_3 inst_cell_123_73 ( BL73, BLN73, WL123);
sram_cell_6t_3 inst_cell_123_72 ( BL72, BLN72, WL123);
sram_cell_6t_3 inst_cell_123_71 ( BL71, BLN71, WL123);
sram_cell_6t_3 inst_cell_123_70 ( BL70, BLN70, WL123);
sram_cell_6t_3 inst_cell_123_69 ( BL69, BLN69, WL123);
sram_cell_6t_3 inst_cell_123_68 ( BL68, BLN68, WL123);
sram_cell_6t_3 inst_cell_123_67 ( BL67, BLN67, WL123);
sram_cell_6t_3 inst_cell_123_66 ( BL66, BLN66, WL123);
sram_cell_6t_3 inst_cell_123_65 ( BL65, BLN65, WL123);
sram_cell_6t_3 inst_cell_123_64 ( BL64, BLN64, WL123);
sram_cell_6t_3 inst_cell_123_63 ( BL63, BLN63, WL123);
sram_cell_6t_3 inst_cell_123_62 ( BL62, BLN62, WL123);
sram_cell_6t_3 inst_cell_123_61 ( BL61, BLN61, WL123);
sram_cell_6t_3 inst_cell_123_60 ( BL60, BLN60, WL123);
sram_cell_6t_3 inst_cell_123_59 ( BL59, BLN59, WL123);
sram_cell_6t_3 inst_cell_123_58 ( BL58, BLN58, WL123);
sram_cell_6t_3 inst_cell_123_57 ( BL57, BLN57, WL123);
sram_cell_6t_3 inst_cell_123_56 ( BL56, BLN56, WL123);
sram_cell_6t_3 inst_cell_123_55 ( BL55, BLN55, WL123);
sram_cell_6t_3 inst_cell_123_54 ( BL54, BLN54, WL123);
sram_cell_6t_3 inst_cell_123_53 ( BL53, BLN53, WL123);
sram_cell_6t_3 inst_cell_123_52 ( BL52, BLN52, WL123);
sram_cell_6t_3 inst_cell_123_51 ( BL51, BLN51, WL123);
sram_cell_6t_3 inst_cell_123_50 ( BL50, BLN50, WL123);
sram_cell_6t_3 inst_cell_123_49 ( BL49, BLN49, WL123);
sram_cell_6t_3 inst_cell_123_48 ( BL48, BLN48, WL123);
sram_cell_6t_3 inst_cell_123_47 ( BL47, BLN47, WL123);
sram_cell_6t_3 inst_cell_123_46 ( BL46, BLN46, WL123);
sram_cell_6t_3 inst_cell_123_45 ( BL45, BLN45, WL123);
sram_cell_6t_3 inst_cell_123_44 ( BL44, BLN44, WL123);
sram_cell_6t_3 inst_cell_123_43 ( BL43, BLN43, WL123);
sram_cell_6t_3 inst_cell_123_42 ( BL42, BLN42, WL123);
sram_cell_6t_3 inst_cell_123_41 ( BL41, BLN41, WL123);
sram_cell_6t_3 inst_cell_123_40 ( BL40, BLN40, WL123);
sram_cell_6t_3 inst_cell_123_39 ( BL39, BLN39, WL123);
sram_cell_6t_3 inst_cell_123_38 ( BL38, BLN38, WL123);
sram_cell_6t_3 inst_cell_123_37 ( BL37, BLN37, WL123);
sram_cell_6t_3 inst_cell_123_36 ( BL36, BLN36, WL123);
sram_cell_6t_3 inst_cell_123_35 ( BL35, BLN35, WL123);
sram_cell_6t_3 inst_cell_123_34 ( BL34, BLN34, WL123);
sram_cell_6t_3 inst_cell_123_33 ( BL33, BLN33, WL123);
sram_cell_6t_3 inst_cell_123_32 ( BL32, BLN32, WL123);
sram_cell_6t_3 inst_cell_123_31 ( BL31, BLN31, WL123);
sram_cell_6t_3 inst_cell_123_30 ( BL30, BLN30, WL123);
sram_cell_6t_3 inst_cell_123_29 ( BL29, BLN29, WL123);
sram_cell_6t_3 inst_cell_123_28 ( BL28, BLN28, WL123);
sram_cell_6t_3 inst_cell_123_27 ( BL27, BLN27, WL123);
sram_cell_6t_3 inst_cell_123_26 ( BL26, BLN26, WL123);
sram_cell_6t_3 inst_cell_123_25 ( BL25, BLN25, WL123);
sram_cell_6t_3 inst_cell_123_24 ( BL24, BLN24, WL123);
sram_cell_6t_3 inst_cell_123_23 ( BL23, BLN23, WL123);
sram_cell_6t_3 inst_cell_123_22 ( BL22, BLN22, WL123);
sram_cell_6t_3 inst_cell_123_21 ( BL21, BLN21, WL123);
sram_cell_6t_3 inst_cell_123_20 ( BL20, BLN20, WL123);
sram_cell_6t_3 inst_cell_123_19 ( BL19, BLN19, WL123);
sram_cell_6t_3 inst_cell_123_18 ( BL18, BLN18, WL123);
sram_cell_6t_3 inst_cell_123_17 ( BL17, BLN17, WL123);
sram_cell_6t_3 inst_cell_123_16 ( BL16, BLN16, WL123);
sram_cell_6t_3 inst_cell_123_15 ( BL15, BLN15, WL123);
sram_cell_6t_3 inst_cell_123_14 ( BL14, BLN14, WL123);
sram_cell_6t_3 inst_cell_123_13 ( BL13, BLN13, WL123);
sram_cell_6t_3 inst_cell_123_12 ( BL12, BLN12, WL123);
sram_cell_6t_3 inst_cell_123_11 ( BL11, BLN11, WL123);
sram_cell_6t_3 inst_cell_123_10 ( BL10, BLN10, WL123);
sram_cell_6t_3 inst_cell_123_9 ( BL9, BLN9, WL123);
sram_cell_6t_3 inst_cell_123_8 ( BL8, BLN8, WL123);
sram_cell_6t_3 inst_cell_123_7 ( BL7, BLN7, WL123);
sram_cell_6t_3 inst_cell_123_6 ( BL6, BLN6, WL123);
sram_cell_6t_3 inst_cell_123_5 ( BL5, BLN5, WL123);
sram_cell_6t_3 inst_cell_123_4 ( BL4, BLN4, WL123);
sram_cell_6t_3 inst_cell_123_3 ( BL3, BLN3, WL123);
sram_cell_6t_3 inst_cell_123_2 ( BL2, BLN2, WL123);
sram_cell_6t_3 inst_cell_123_1 ( BL1, BLN1, WL123);
sram_cell_6t_3 inst_cell_123_0 ( BL0, BLN0, WL123);
sram_cell_6t_3 inst_cell_122_127 ( BL127, BLN127, WL122);
sram_cell_6t_3 inst_cell_122_126 ( BL126, BLN126, WL122);
sram_cell_6t_3 inst_cell_122_125 ( BL125, BLN125, WL122);
sram_cell_6t_3 inst_cell_122_124 ( BL124, BLN124, WL122);
sram_cell_6t_3 inst_cell_122_123 ( BL123, BLN123, WL122);
sram_cell_6t_3 inst_cell_122_122 ( BL122, BLN122, WL122);
sram_cell_6t_3 inst_cell_122_121 ( BL121, BLN121, WL122);
sram_cell_6t_3 inst_cell_122_120 ( BL120, BLN120, WL122);
sram_cell_6t_3 inst_cell_122_119 ( BL119, BLN119, WL122);
sram_cell_6t_3 inst_cell_122_118 ( BL118, BLN118, WL122);
sram_cell_6t_3 inst_cell_122_117 ( BL117, BLN117, WL122);
sram_cell_6t_3 inst_cell_122_116 ( BL116, BLN116, WL122);
sram_cell_6t_3 inst_cell_122_115 ( BL115, BLN115, WL122);
sram_cell_6t_3 inst_cell_122_114 ( BL114, BLN114, WL122);
sram_cell_6t_3 inst_cell_122_113 ( BL113, BLN113, WL122);
sram_cell_6t_3 inst_cell_122_112 ( BL112, BLN112, WL122);
sram_cell_6t_3 inst_cell_122_111 ( BL111, BLN111, WL122);
sram_cell_6t_3 inst_cell_122_110 ( BL110, BLN110, WL122);
sram_cell_6t_3 inst_cell_122_109 ( BL109, BLN109, WL122);
sram_cell_6t_3 inst_cell_122_108 ( BL108, BLN108, WL122);
sram_cell_6t_3 inst_cell_122_107 ( BL107, BLN107, WL122);
sram_cell_6t_3 inst_cell_122_106 ( BL106, BLN106, WL122);
sram_cell_6t_3 inst_cell_122_105 ( BL105, BLN105, WL122);
sram_cell_6t_3 inst_cell_122_104 ( BL104, BLN104, WL122);
sram_cell_6t_3 inst_cell_122_103 ( BL103, BLN103, WL122);
sram_cell_6t_3 inst_cell_122_102 ( BL102, BLN102, WL122);
sram_cell_6t_3 inst_cell_122_101 ( BL101, BLN101, WL122);
sram_cell_6t_3 inst_cell_122_100 ( BL100, BLN100, WL122);
sram_cell_6t_3 inst_cell_122_99 ( BL99, BLN99, WL122);
sram_cell_6t_3 inst_cell_122_98 ( BL98, BLN98, WL122);
sram_cell_6t_3 inst_cell_122_97 ( BL97, BLN97, WL122);
sram_cell_6t_3 inst_cell_122_96 ( BL96, BLN96, WL122);
sram_cell_6t_3 inst_cell_122_95 ( BL95, BLN95, WL122);
sram_cell_6t_3 inst_cell_122_94 ( BL94, BLN94, WL122);
sram_cell_6t_3 inst_cell_122_93 ( BL93, BLN93, WL122);
sram_cell_6t_3 inst_cell_122_92 ( BL92, BLN92, WL122);
sram_cell_6t_3 inst_cell_122_91 ( BL91, BLN91, WL122);
sram_cell_6t_3 inst_cell_122_90 ( BL90, BLN90, WL122);
sram_cell_6t_3 inst_cell_122_89 ( BL89, BLN89, WL122);
sram_cell_6t_3 inst_cell_122_88 ( BL88, BLN88, WL122);
sram_cell_6t_3 inst_cell_122_87 ( BL87, BLN87, WL122);
sram_cell_6t_3 inst_cell_122_86 ( BL86, BLN86, WL122);
sram_cell_6t_3 inst_cell_122_85 ( BL85, BLN85, WL122);
sram_cell_6t_3 inst_cell_122_84 ( BL84, BLN84, WL122);
sram_cell_6t_3 inst_cell_122_83 ( BL83, BLN83, WL122);
sram_cell_6t_3 inst_cell_122_82 ( BL82, BLN82, WL122);
sram_cell_6t_3 inst_cell_122_81 ( BL81, BLN81, WL122);
sram_cell_6t_3 inst_cell_122_80 ( BL80, BLN80, WL122);
sram_cell_6t_3 inst_cell_122_79 ( BL79, BLN79, WL122);
sram_cell_6t_3 inst_cell_122_78 ( BL78, BLN78, WL122);
sram_cell_6t_3 inst_cell_122_77 ( BL77, BLN77, WL122);
sram_cell_6t_3 inst_cell_122_76 ( BL76, BLN76, WL122);
sram_cell_6t_3 inst_cell_122_75 ( BL75, BLN75, WL122);
sram_cell_6t_3 inst_cell_122_74 ( BL74, BLN74, WL122);
sram_cell_6t_3 inst_cell_122_73 ( BL73, BLN73, WL122);
sram_cell_6t_3 inst_cell_122_72 ( BL72, BLN72, WL122);
sram_cell_6t_3 inst_cell_122_71 ( BL71, BLN71, WL122);
sram_cell_6t_3 inst_cell_122_70 ( BL70, BLN70, WL122);
sram_cell_6t_3 inst_cell_122_69 ( BL69, BLN69, WL122);
sram_cell_6t_3 inst_cell_122_68 ( BL68, BLN68, WL122);
sram_cell_6t_3 inst_cell_122_67 ( BL67, BLN67, WL122);
sram_cell_6t_3 inst_cell_122_66 ( BL66, BLN66, WL122);
sram_cell_6t_3 inst_cell_122_65 ( BL65, BLN65, WL122);
sram_cell_6t_3 inst_cell_122_64 ( BL64, BLN64, WL122);
sram_cell_6t_3 inst_cell_122_63 ( BL63, BLN63, WL122);
sram_cell_6t_3 inst_cell_122_62 ( BL62, BLN62, WL122);
sram_cell_6t_3 inst_cell_122_61 ( BL61, BLN61, WL122);
sram_cell_6t_3 inst_cell_122_60 ( BL60, BLN60, WL122);
sram_cell_6t_3 inst_cell_122_59 ( BL59, BLN59, WL122);
sram_cell_6t_3 inst_cell_122_58 ( BL58, BLN58, WL122);
sram_cell_6t_3 inst_cell_122_57 ( BL57, BLN57, WL122);
sram_cell_6t_3 inst_cell_122_56 ( BL56, BLN56, WL122);
sram_cell_6t_3 inst_cell_122_55 ( BL55, BLN55, WL122);
sram_cell_6t_3 inst_cell_122_54 ( BL54, BLN54, WL122);
sram_cell_6t_3 inst_cell_122_53 ( BL53, BLN53, WL122);
sram_cell_6t_3 inst_cell_122_52 ( BL52, BLN52, WL122);
sram_cell_6t_3 inst_cell_122_51 ( BL51, BLN51, WL122);
sram_cell_6t_3 inst_cell_122_50 ( BL50, BLN50, WL122);
sram_cell_6t_3 inst_cell_122_49 ( BL49, BLN49, WL122);
sram_cell_6t_3 inst_cell_122_48 ( BL48, BLN48, WL122);
sram_cell_6t_3 inst_cell_127_3 ( BL3, BLN3, WL127);
sram_cell_6t_3 inst_cell_122_3 ( BL3, BLN3, WL122);
sram_cell_6t_3 inst_cell_127_2 ( BL2, BLN2, WL127);
sram_cell_6t_3 inst_cell_122_2 ( BL2, BLN2, WL122);
sram_cell_6t_3 inst_cell_127_1 ( BL1, BLN1, WL127);
sram_cell_6t_3 inst_cell_122_1 ( BL1, BLN1, WL122);
sram_cell_6t_3 inst_cell_127_0 ( BL0, BLN0, WL127);
sram_cell_6t_3 inst_cell_122_0 ( BL0, BLN0, WL122);
sram_cell_6t_3 inst_cell_122_47 ( BL47, BLN47, WL122);
sram_cell_6t_3 inst_cell_122_46 ( BL46, BLN46, WL122);
sram_cell_6t_3 inst_cell_122_45 ( BL45, BLN45, WL122);
sram_cell_6t_3 inst_cell_122_44 ( BL44, BLN44, WL122);
sram_cell_6t_3 inst_cell_122_43 ( BL43, BLN43, WL122);
sram_cell_6t_3 inst_cell_122_42 ( BL42, BLN42, WL122);
sram_cell_6t_3 inst_cell_122_41 ( BL41, BLN41, WL122);
sram_cell_6t_3 inst_cell_122_40 ( BL40, BLN40, WL122);
sram_cell_6t_3 inst_cell_122_39 ( BL39, BLN39, WL122);
sram_cell_6t_3 inst_cell_122_38 ( BL38, BLN38, WL122);
sram_cell_6t_3 inst_cell_122_37 ( BL37, BLN37, WL122);
sram_cell_6t_3 inst_cell_122_36 ( BL36, BLN36, WL122);
sram_cell_6t_3 inst_cell_122_35 ( BL35, BLN35, WL122);
sram_cell_6t_3 inst_cell_122_34 ( BL34, BLN34, WL122);
sram_cell_6t_3 inst_cell_122_33 ( BL33, BLN33, WL122);
sram_cell_6t_3 inst_cell_122_32 ( BL32, BLN32, WL122);
sram_cell_6t_3 inst_cell_122_31 ( BL31, BLN31, WL122);
sram_cell_6t_3 inst_cell_122_30 ( BL30, BLN30, WL122);
sram_cell_6t_3 inst_cell_122_29 ( BL29, BLN29, WL122);
sram_cell_6t_3 inst_cell_122_28 ( BL28, BLN28, WL122);
sram_cell_6t_3 inst_cell_122_27 ( BL27, BLN27, WL122);
sram_cell_6t_3 inst_cell_122_26 ( BL26, BLN26, WL122);
sram_cell_6t_3 inst_cell_122_25 ( BL25, BLN25, WL122);
sram_cell_6t_3 inst_cell_122_24 ( BL24, BLN24, WL122);
sram_cell_6t_3 inst_cell_122_23 ( BL23, BLN23, WL122);
sram_cell_6t_3 inst_cell_122_22 ( BL22, BLN22, WL122);
sram_cell_6t_3 inst_cell_122_21 ( BL21, BLN21, WL122);
sram_cell_6t_3 inst_cell_122_20 ( BL20, BLN20, WL122);
sram_cell_6t_3 inst_cell_122_19 ( BL19, BLN19, WL122);
sram_cell_6t_3 inst_cell_122_18 ( BL18, BLN18, WL122);
sram_cell_6t_3 inst_cell_122_17 ( BL17, BLN17, WL122);
sram_cell_6t_3 inst_cell_122_16 ( BL16, BLN16, WL122);
sram_cell_6t_3 inst_cell_122_15 ( BL15, BLN15, WL122);
sram_cell_6t_3 inst_cell_122_14 ( BL14, BLN14, WL122);
sram_cell_6t_3 inst_cell_122_13 ( BL13, BLN13, WL122);
sram_cell_6t_3 inst_cell_122_12 ( BL12, BLN12, WL122);
sram_cell_6t_3 inst_cell_122_11 ( BL11, BLN11, WL122);
sram_cell_6t_3 inst_cell_122_10 ( BL10, BLN10, WL122);
sram_cell_6t_3 inst_cell_122_9 ( BL9, BLN9, WL122);
sram_cell_6t_3 inst_cell_122_8 ( BL8, BLN8, WL122);
sram_cell_6t_3 inst_cell_122_7 ( BL7, BLN7, WL122);
sram_cell_6t_3 inst_cell_122_6 ( BL6, BLN6, WL122);
sram_cell_6t_3 inst_cell_122_5 ( BL5, BLN5, WL122);
sram_cell_6t_3 inst_cell_122_4 ( BL4, BLN4, WL122);
sram_cell_6t_3 inst_cell_121_127 ( BL127, BLN127, WL121);
sram_cell_6t_3 inst_cell_121_126 ( BL126, BLN126, WL121);
sram_cell_6t_3 inst_cell_121_125 ( BL125, BLN125, WL121);
sram_cell_6t_3 inst_cell_121_124 ( BL124, BLN124, WL121);
sram_cell_6t_3 inst_cell_121_123 ( BL123, BLN123, WL121);
sram_cell_6t_3 inst_cell_121_122 ( BL122, BLN122, WL121);
sram_cell_6t_3 inst_cell_121_121 ( BL121, BLN121, WL121);
sram_cell_6t_3 inst_cell_121_120 ( BL120, BLN120, WL121);
sram_cell_6t_3 inst_cell_121_119 ( BL119, BLN119, WL121);
sram_cell_6t_3 inst_cell_121_118 ( BL118, BLN118, WL121);
sram_cell_6t_3 inst_cell_121_117 ( BL117, BLN117, WL121);
sram_cell_6t_3 inst_cell_121_116 ( BL116, BLN116, WL121);
sram_cell_6t_3 inst_cell_121_115 ( BL115, BLN115, WL121);
sram_cell_6t_3 inst_cell_121_114 ( BL114, BLN114, WL121);
sram_cell_6t_3 inst_cell_121_113 ( BL113, BLN113, WL121);
sram_cell_6t_3 inst_cell_121_112 ( BL112, BLN112, WL121);
sram_cell_6t_3 inst_cell_121_111 ( BL111, BLN111, WL121);
sram_cell_6t_3 inst_cell_121_110 ( BL110, BLN110, WL121);
sram_cell_6t_3 inst_cell_121_109 ( BL109, BLN109, WL121);
sram_cell_6t_3 inst_cell_121_108 ( BL108, BLN108, WL121);
sram_cell_6t_3 inst_cell_121_107 ( BL107, BLN107, WL121);
sram_cell_6t_3 inst_cell_121_106 ( BL106, BLN106, WL121);
sram_cell_6t_3 inst_cell_121_105 ( BL105, BLN105, WL121);
sram_cell_6t_3 inst_cell_121_104 ( BL104, BLN104, WL121);
sram_cell_6t_3 inst_cell_121_103 ( BL103, BLN103, WL121);
sram_cell_6t_3 inst_cell_121_102 ( BL102, BLN102, WL121);
sram_cell_6t_3 inst_cell_121_101 ( BL101, BLN101, WL121);
sram_cell_6t_3 inst_cell_121_100 ( BL100, BLN100, WL121);
sram_cell_6t_3 inst_cell_121_99 ( BL99, BLN99, WL121);
sram_cell_6t_3 inst_cell_121_98 ( BL98, BLN98, WL121);
sram_cell_6t_3 inst_cell_121_97 ( BL97, BLN97, WL121);
sram_cell_6t_3 inst_cell_121_96 ( BL96, BLN96, WL121);
sram_cell_6t_3 inst_cell_121_95 ( BL95, BLN95, WL121);
sram_cell_6t_3 inst_cell_121_94 ( BL94, BLN94, WL121);
sram_cell_6t_3 inst_cell_121_93 ( BL93, BLN93, WL121);
sram_cell_6t_3 inst_cell_121_92 ( BL92, BLN92, WL121);
sram_cell_6t_3 inst_cell_121_91 ( BL91, BLN91, WL121);
sram_cell_6t_3 inst_cell_121_90 ( BL90, BLN90, WL121);
sram_cell_6t_3 inst_cell_121_89 ( BL89, BLN89, WL121);
sram_cell_6t_3 inst_cell_121_88 ( BL88, BLN88, WL121);
sram_cell_6t_3 inst_cell_121_87 ( BL87, BLN87, WL121);
sram_cell_6t_3 inst_cell_121_86 ( BL86, BLN86, WL121);
sram_cell_6t_3 inst_cell_121_85 ( BL85, BLN85, WL121);
sram_cell_6t_3 inst_cell_121_84 ( BL84, BLN84, WL121);
sram_cell_6t_3 inst_cell_121_83 ( BL83, BLN83, WL121);
sram_cell_6t_3 inst_cell_121_82 ( BL82, BLN82, WL121);
sram_cell_6t_3 inst_cell_121_81 ( BL81, BLN81, WL121);
sram_cell_6t_3 inst_cell_121_80 ( BL80, BLN80, WL121);
sram_cell_6t_3 inst_cell_121_79 ( BL79, BLN79, WL121);
sram_cell_6t_3 inst_cell_121_78 ( BL78, BLN78, WL121);
sram_cell_6t_3 inst_cell_121_77 ( BL77, BLN77, WL121);
sram_cell_6t_3 inst_cell_121_76 ( BL76, BLN76, WL121);
sram_cell_6t_3 inst_cell_121_75 ( BL75, BLN75, WL121);
sram_cell_6t_3 inst_cell_121_74 ( BL74, BLN74, WL121);
sram_cell_6t_3 inst_cell_121_73 ( BL73, BLN73, WL121);
sram_cell_6t_3 inst_cell_121_72 ( BL72, BLN72, WL121);
sram_cell_6t_3 inst_cell_121_71 ( BL71, BLN71, WL121);
sram_cell_6t_3 inst_cell_121_70 ( BL70, BLN70, WL121);
sram_cell_6t_3 inst_cell_121_69 ( BL69, BLN69, WL121);
sram_cell_6t_3 inst_cell_121_68 ( BL68, BLN68, WL121);
sram_cell_6t_3 inst_cell_121_67 ( BL67, BLN67, WL121);
sram_cell_6t_3 inst_cell_121_66 ( BL66, BLN66, WL121);
sram_cell_6t_3 inst_cell_121_65 ( BL65, BLN65, WL121);
sram_cell_6t_3 inst_cell_121_64 ( BL64, BLN64, WL121);
sram_cell_6t_3 inst_cell_121_63 ( BL63, BLN63, WL121);
sram_cell_6t_3 inst_cell_121_62 ( BL62, BLN62, WL121);
sram_cell_6t_3 inst_cell_121_61 ( BL61, BLN61, WL121);
sram_cell_6t_3 inst_cell_121_60 ( BL60, BLN60, WL121);
sram_cell_6t_3 inst_cell_121_59 ( BL59, BLN59, WL121);
sram_cell_6t_3 inst_cell_121_58 ( BL58, BLN58, WL121);
sram_cell_6t_3 inst_cell_121_57 ( BL57, BLN57, WL121);
sram_cell_6t_3 inst_cell_121_56 ( BL56, BLN56, WL121);
sram_cell_6t_3 inst_cell_121_55 ( BL55, BLN55, WL121);
sram_cell_6t_3 inst_cell_121_54 ( BL54, BLN54, WL121);
sram_cell_6t_3 inst_cell_121_53 ( BL53, BLN53, WL121);
sram_cell_6t_3 inst_cell_121_52 ( BL52, BLN52, WL121);
sram_cell_6t_3 inst_cell_121_51 ( BL51, BLN51, WL121);
sram_cell_6t_3 inst_cell_121_50 ( BL50, BLN50, WL121);
sram_cell_6t_3 inst_cell_121_49 ( BL49, BLN49, WL121);
sram_cell_6t_3 inst_cell_121_48 ( BL48, BLN48, WL121);
sram_cell_6t_3 inst_cell_121_47 ( BL47, BLN47, WL121);
sram_cell_6t_3 inst_cell_121_46 ( BL46, BLN46, WL121);
sram_cell_6t_3 inst_cell_121_45 ( BL45, BLN45, WL121);
sram_cell_6t_3 inst_cell_121_44 ( BL44, BLN44, WL121);
sram_cell_6t_3 inst_cell_121_43 ( BL43, BLN43, WL121);
sram_cell_6t_3 inst_cell_121_42 ( BL42, BLN42, WL121);
sram_cell_6t_3 inst_cell_121_41 ( BL41, BLN41, WL121);
sram_cell_6t_3 inst_cell_121_40 ( BL40, BLN40, WL121);
sram_cell_6t_3 inst_cell_121_39 ( BL39, BLN39, WL121);
sram_cell_6t_3 inst_cell_121_38 ( BL38, BLN38, WL121);
sram_cell_6t_3 inst_cell_121_37 ( BL37, BLN37, WL121);
sram_cell_6t_3 inst_cell_121_36 ( BL36, BLN36, WL121);
sram_cell_6t_3 inst_cell_121_35 ( BL35, BLN35, WL121);
sram_cell_6t_3 inst_cell_121_34 ( BL34, BLN34, WL121);
sram_cell_6t_3 inst_cell_121_33 ( BL33, BLN33, WL121);
sram_cell_6t_3 inst_cell_121_32 ( BL32, BLN32, WL121);
sram_cell_6t_3 inst_cell_121_31 ( BL31, BLN31, WL121);
sram_cell_6t_3 inst_cell_121_30 ( BL30, BLN30, WL121);
sram_cell_6t_3 inst_cell_121_29 ( BL29, BLN29, WL121);
sram_cell_6t_3 inst_cell_121_28 ( BL28, BLN28, WL121);
sram_cell_6t_3 inst_cell_121_27 ( BL27, BLN27, WL121);
sram_cell_6t_3 inst_cell_121_26 ( BL26, BLN26, WL121);
sram_cell_6t_3 inst_cell_121_25 ( BL25, BLN25, WL121);
sram_cell_6t_3 inst_cell_121_24 ( BL24, BLN24, WL121);
sram_cell_6t_3 inst_cell_121_23 ( BL23, BLN23, WL121);
sram_cell_6t_3 inst_cell_121_22 ( BL22, BLN22, WL121);
sram_cell_6t_3 inst_cell_121_21 ( BL21, BLN21, WL121);
sram_cell_6t_3 inst_cell_121_20 ( BL20, BLN20, WL121);
sram_cell_6t_3 inst_cell_121_19 ( BL19, BLN19, WL121);
sram_cell_6t_3 inst_cell_121_18 ( BL18, BLN18, WL121);
sram_cell_6t_3 inst_cell_121_17 ( BL17, BLN17, WL121);
sram_cell_6t_3 inst_cell_121_16 ( BL16, BLN16, WL121);
sram_cell_6t_3 inst_cell_121_15 ( BL15, BLN15, WL121);
sram_cell_6t_3 inst_cell_121_14 ( BL14, BLN14, WL121);
sram_cell_6t_3 inst_cell_121_13 ( BL13, BLN13, WL121);
sram_cell_6t_3 inst_cell_121_12 ( BL12, BLN12, WL121);
sram_cell_6t_3 inst_cell_121_11 ( BL11, BLN11, WL121);
sram_cell_6t_3 inst_cell_121_10 ( BL10, BLN10, WL121);
sram_cell_6t_3 inst_cell_121_9 ( BL9, BLN9, WL121);
sram_cell_6t_3 inst_cell_121_8 ( BL8, BLN8, WL121);
sram_cell_6t_3 inst_cell_121_7 ( BL7, BLN7, WL121);
sram_cell_6t_3 inst_cell_121_6 ( BL6, BLN6, WL121);
sram_cell_6t_3 inst_cell_121_5 ( BL5, BLN5, WL121);
sram_cell_6t_3 inst_cell_121_4 ( BL4, BLN4, WL121);
sram_cell_6t_3 inst_cell_121_3 ( BL3, BLN3, WL121);
sram_cell_6t_3 inst_cell_121_2 ( BL2, BLN2, WL121);
sram_cell_6t_3 inst_cell_121_1 ( BL1, BLN1, WL121);
sram_cell_6t_3 inst_cell_121_0 ( BL0, BLN0, WL121);
sram_cell_6t_3 inst_cell_120_127 ( BL127, BLN127, WL120);
sram_cell_6t_3 inst_cell_120_126 ( BL126, BLN126, WL120);
sram_cell_6t_3 inst_cell_120_125 ( BL125, BLN125, WL120);
sram_cell_6t_3 inst_cell_120_124 ( BL124, BLN124, WL120);
sram_cell_6t_3 inst_cell_120_123 ( BL123, BLN123, WL120);
sram_cell_6t_3 inst_cell_120_122 ( BL122, BLN122, WL120);
sram_cell_6t_3 inst_cell_120_121 ( BL121, BLN121, WL120);
sram_cell_6t_3 inst_cell_120_120 ( BL120, BLN120, WL120);
sram_cell_6t_3 inst_cell_120_119 ( BL119, BLN119, WL120);
sram_cell_6t_3 inst_cell_120_118 ( BL118, BLN118, WL120);
sram_cell_6t_3 inst_cell_120_117 ( BL117, BLN117, WL120);
sram_cell_6t_3 inst_cell_120_116 ( BL116, BLN116, WL120);
sram_cell_6t_3 inst_cell_120_115 ( BL115, BLN115, WL120);
sram_cell_6t_3 inst_cell_120_114 ( BL114, BLN114, WL120);
sram_cell_6t_3 inst_cell_120_113 ( BL113, BLN113, WL120);
sram_cell_6t_3 inst_cell_120_112 ( BL112, BLN112, WL120);
sram_cell_6t_3 inst_cell_120_111 ( BL111, BLN111, WL120);
sram_cell_6t_3 inst_cell_120_110 ( BL110, BLN110, WL120);
sram_cell_6t_3 inst_cell_120_109 ( BL109, BLN109, WL120);
sram_cell_6t_3 inst_cell_120_108 ( BL108, BLN108, WL120);
sram_cell_6t_3 inst_cell_120_107 ( BL107, BLN107, WL120);
sram_cell_6t_3 inst_cell_120_106 ( BL106, BLN106, WL120);
sram_cell_6t_3 inst_cell_120_105 ( BL105, BLN105, WL120);
sram_cell_6t_3 inst_cell_120_104 ( BL104, BLN104, WL120);
sram_cell_6t_3 inst_cell_120_103 ( BL103, BLN103, WL120);
sram_cell_6t_3 inst_cell_120_102 ( BL102, BLN102, WL120);
sram_cell_6t_3 inst_cell_120_101 ( BL101, BLN101, WL120);
sram_cell_6t_3 inst_cell_120_100 ( BL100, BLN100, WL120);
sram_cell_6t_3 inst_cell_120_99 ( BL99, BLN99, WL120);
sram_cell_6t_3 inst_cell_120_98 ( BL98, BLN98, WL120);
sram_cell_6t_3 inst_cell_120_97 ( BL97, BLN97, WL120);
sram_cell_6t_3 inst_cell_120_96 ( BL96, BLN96, WL120);
sram_cell_6t_3 inst_cell_120_95 ( BL95, BLN95, WL120);
sram_cell_6t_3 inst_cell_120_94 ( BL94, BLN94, WL120);
sram_cell_6t_3 inst_cell_120_93 ( BL93, BLN93, WL120);
sram_cell_6t_3 inst_cell_120_92 ( BL92, BLN92, WL120);
sram_cell_6t_3 inst_cell_120_91 ( BL91, BLN91, WL120);
sram_cell_6t_3 inst_cell_120_90 ( BL90, BLN90, WL120);
sram_cell_6t_3 inst_cell_120_89 ( BL89, BLN89, WL120);
sram_cell_6t_3 inst_cell_120_88 ( BL88, BLN88, WL120);
sram_cell_6t_3 inst_cell_120_87 ( BL87, BLN87, WL120);
sram_cell_6t_3 inst_cell_120_86 ( BL86, BLN86, WL120);
sram_cell_6t_3 inst_cell_120_85 ( BL85, BLN85, WL120);
sram_cell_6t_3 inst_cell_120_84 ( BL84, BLN84, WL120);
sram_cell_6t_3 inst_cell_120_83 ( BL83, BLN83, WL120);
sram_cell_6t_3 inst_cell_120_82 ( BL82, BLN82, WL120);
sram_cell_6t_3 inst_cell_120_81 ( BL81, BLN81, WL120);
sram_cell_6t_3 inst_cell_120_80 ( BL80, BLN80, WL120);
sram_cell_6t_3 inst_cell_120_79 ( BL79, BLN79, WL120);
sram_cell_6t_3 inst_cell_120_78 ( BL78, BLN78, WL120);
sram_cell_6t_3 inst_cell_120_77 ( BL77, BLN77, WL120);
sram_cell_6t_3 inst_cell_120_76 ( BL76, BLN76, WL120);
sram_cell_6t_3 inst_cell_120_75 ( BL75, BLN75, WL120);
sram_cell_6t_3 inst_cell_120_74 ( BL74, BLN74, WL120);
sram_cell_6t_3 inst_cell_120_73 ( BL73, BLN73, WL120);
sram_cell_6t_3 inst_cell_120_72 ( BL72, BLN72, WL120);
sram_cell_6t_3 inst_cell_120_71 ( BL71, BLN71, WL120);
sram_cell_6t_3 inst_cell_120_70 ( BL70, BLN70, WL120);
sram_cell_6t_3 inst_cell_120_69 ( BL69, BLN69, WL120);
sram_cell_6t_3 inst_cell_120_68 ( BL68, BLN68, WL120);
sram_cell_6t_3 inst_cell_120_67 ( BL67, BLN67, WL120);
sram_cell_6t_3 inst_cell_120_66 ( BL66, BLN66, WL120);
sram_cell_6t_3 inst_cell_120_65 ( BL65, BLN65, WL120);
sram_cell_6t_3 inst_cell_120_64 ( BL64, BLN64, WL120);
sram_cell_6t_3 inst_cell_120_63 ( BL63, BLN63, WL120);
sram_cell_6t_3 inst_cell_120_62 ( BL62, BLN62, WL120);
sram_cell_6t_3 inst_cell_120_61 ( BL61, BLN61, WL120);
sram_cell_6t_3 inst_cell_120_60 ( BL60, BLN60, WL120);
sram_cell_6t_3 inst_cell_120_59 ( BL59, BLN59, WL120);
sram_cell_6t_3 inst_cell_120_58 ( BL58, BLN58, WL120);
sram_cell_6t_3 inst_cell_120_57 ( BL57, BLN57, WL120);
sram_cell_6t_3 inst_cell_120_56 ( BL56, BLN56, WL120);
sram_cell_6t_3 inst_cell_120_55 ( BL55, BLN55, WL120);
sram_cell_6t_3 inst_cell_120_54 ( BL54, BLN54, WL120);
sram_cell_6t_3 inst_cell_120_53 ( BL53, BLN53, WL120);
sram_cell_6t_3 inst_cell_120_52 ( BL52, BLN52, WL120);
sram_cell_6t_3 inst_cell_120_51 ( BL51, BLN51, WL120);
sram_cell_6t_3 inst_cell_120_50 ( BL50, BLN50, WL120);
sram_cell_6t_3 inst_cell_120_49 ( BL49, BLN49, WL120);
sram_cell_6t_3 inst_cell_120_48 ( BL48, BLN48, WL120);
sram_cell_6t_3 inst_cell_120_47 ( BL47, BLN47, WL120);
sram_cell_6t_3 inst_cell_120_46 ( BL46, BLN46, WL120);
sram_cell_6t_3 inst_cell_120_45 ( BL45, BLN45, WL120);
sram_cell_6t_3 inst_cell_120_44 ( BL44, BLN44, WL120);
sram_cell_6t_3 inst_cell_120_43 ( BL43, BLN43, WL120);
sram_cell_6t_3 inst_cell_120_42 ( BL42, BLN42, WL120);
sram_cell_6t_3 inst_cell_120_41 ( BL41, BLN41, WL120);
sram_cell_6t_3 inst_cell_120_40 ( BL40, BLN40, WL120);
sram_cell_6t_3 inst_cell_120_39 ( BL39, BLN39, WL120);
sram_cell_6t_3 inst_cell_120_38 ( BL38, BLN38, WL120);
sram_cell_6t_3 inst_cell_120_37 ( BL37, BLN37, WL120);
sram_cell_6t_3 inst_cell_120_36 ( BL36, BLN36, WL120);
sram_cell_6t_3 inst_cell_120_35 ( BL35, BLN35, WL120);
sram_cell_6t_3 inst_cell_120_34 ( BL34, BLN34, WL120);
sram_cell_6t_3 inst_cell_120_33 ( BL33, BLN33, WL120);
sram_cell_6t_3 inst_cell_120_32 ( BL32, BLN32, WL120);
sram_cell_6t_3 inst_cell_120_31 ( BL31, BLN31, WL120);
sram_cell_6t_3 inst_cell_120_30 ( BL30, BLN30, WL120);
sram_cell_6t_3 inst_cell_120_29 ( BL29, BLN29, WL120);
sram_cell_6t_3 inst_cell_120_28 ( BL28, BLN28, WL120);
sram_cell_6t_3 inst_cell_120_27 ( BL27, BLN27, WL120);
sram_cell_6t_3 inst_cell_120_26 ( BL26, BLN26, WL120);
sram_cell_6t_3 inst_cell_120_25 ( BL25, BLN25, WL120);
sram_cell_6t_3 inst_cell_120_24 ( BL24, BLN24, WL120);
sram_cell_6t_3 inst_cell_120_23 ( BL23, BLN23, WL120);
sram_cell_6t_3 inst_cell_120_22 ( BL22, BLN22, WL120);
sram_cell_6t_3 inst_cell_120_21 ( BL21, BLN21, WL120);
sram_cell_6t_3 inst_cell_120_20 ( BL20, BLN20, WL120);
sram_cell_6t_3 inst_cell_120_19 ( BL19, BLN19, WL120);
sram_cell_6t_3 inst_cell_120_18 ( BL18, BLN18, WL120);
sram_cell_6t_3 inst_cell_120_17 ( BL17, BLN17, WL120);
sram_cell_6t_3 inst_cell_120_16 ( BL16, BLN16, WL120);
sram_cell_6t_3 inst_cell_120_15 ( BL15, BLN15, WL120);
sram_cell_6t_3 inst_cell_120_14 ( BL14, BLN14, WL120);
sram_cell_6t_3 inst_cell_120_13 ( BL13, BLN13, WL120);
sram_cell_6t_3 inst_cell_120_12 ( BL12, BLN12, WL120);
sram_cell_6t_3 inst_cell_120_11 ( BL11, BLN11, WL120);
sram_cell_6t_3 inst_cell_120_10 ( BL10, BLN10, WL120);
sram_cell_6t_3 inst_cell_120_9 ( BL9, BLN9, WL120);
sram_cell_6t_3 inst_cell_120_8 ( BL8, BLN8, WL120);
sram_cell_6t_3 inst_cell_120_7 ( BL7, BLN7, WL120);
sram_cell_6t_3 inst_cell_120_6 ( BL6, BLN6, WL120);
sram_cell_6t_3 inst_cell_120_5 ( BL5, BLN5, WL120);
sram_cell_6t_3 inst_cell_120_4 ( BL4, BLN4, WL120);
sram_cell_6t_3 inst_cell_120_3 ( BL3, BLN3, WL120);
sram_cell_6t_3 inst_cell_120_2 ( BL2, BLN2, WL120);
sram_cell_6t_3 inst_cell_120_1 ( BL1, BLN1, WL120);
sram_cell_6t_3 inst_cell_120_0 ( BL0, BLN0, WL120);
sram_cell_6t_3 inst_cell_119_127 ( BL127, BLN127, WL119);
sram_cell_6t_3 inst_cell_119_126 ( BL126, BLN126, WL119);
sram_cell_6t_3 inst_cell_119_125 ( BL125, BLN125, WL119);
sram_cell_6t_3 inst_cell_119_124 ( BL124, BLN124, WL119);
sram_cell_6t_3 inst_cell_119_123 ( BL123, BLN123, WL119);
sram_cell_6t_3 inst_cell_119_122 ( BL122, BLN122, WL119);
sram_cell_6t_3 inst_cell_119_121 ( BL121, BLN121, WL119);
sram_cell_6t_3 inst_cell_119_120 ( BL120, BLN120, WL119);
sram_cell_6t_3 inst_cell_119_119 ( BL119, BLN119, WL119);
sram_cell_6t_3 inst_cell_119_118 ( BL118, BLN118, WL119);
sram_cell_6t_3 inst_cell_119_117 ( BL117, BLN117, WL119);
sram_cell_6t_3 inst_cell_119_116 ( BL116, BLN116, WL119);
sram_cell_6t_3 inst_cell_119_115 ( BL115, BLN115, WL119);
sram_cell_6t_3 inst_cell_119_114 ( BL114, BLN114, WL119);
sram_cell_6t_3 inst_cell_119_113 ( BL113, BLN113, WL119);
sram_cell_6t_3 inst_cell_119_112 ( BL112, BLN112, WL119);
sram_cell_6t_3 inst_cell_119_111 ( BL111, BLN111, WL119);
sram_cell_6t_3 inst_cell_119_110 ( BL110, BLN110, WL119);
sram_cell_6t_3 inst_cell_119_109 ( BL109, BLN109, WL119);
sram_cell_6t_3 inst_cell_119_108 ( BL108, BLN108, WL119);
sram_cell_6t_3 inst_cell_119_107 ( BL107, BLN107, WL119);
sram_cell_6t_3 inst_cell_119_106 ( BL106, BLN106, WL119);
sram_cell_6t_3 inst_cell_119_105 ( BL105, BLN105, WL119);
sram_cell_6t_3 inst_cell_119_104 ( BL104, BLN104, WL119);
sram_cell_6t_3 inst_cell_119_103 ( BL103, BLN103, WL119);
sram_cell_6t_3 inst_cell_119_102 ( BL102, BLN102, WL119);
sram_cell_6t_3 inst_cell_119_101 ( BL101, BLN101, WL119);
sram_cell_6t_3 inst_cell_119_100 ( BL100, BLN100, WL119);
sram_cell_6t_3 inst_cell_119_99 ( BL99, BLN99, WL119);
sram_cell_6t_3 inst_cell_119_98 ( BL98, BLN98, WL119);
sram_cell_6t_3 inst_cell_119_97 ( BL97, BLN97, WL119);
sram_cell_6t_3 inst_cell_119_96 ( BL96, BLN96, WL119);
sram_cell_6t_3 inst_cell_119_95 ( BL95, BLN95, WL119);
sram_cell_6t_3 inst_cell_119_94 ( BL94, BLN94, WL119);
sram_cell_6t_3 inst_cell_119_93 ( BL93, BLN93, WL119);
sram_cell_6t_3 inst_cell_119_92 ( BL92, BLN92, WL119);
sram_cell_6t_3 inst_cell_119_91 ( BL91, BLN91, WL119);
sram_cell_6t_3 inst_cell_119_90 ( BL90, BLN90, WL119);
sram_cell_6t_3 inst_cell_119_89 ( BL89, BLN89, WL119);
sram_cell_6t_3 inst_cell_119_88 ( BL88, BLN88, WL119);
sram_cell_6t_3 inst_cell_119_87 ( BL87, BLN87, WL119);
sram_cell_6t_3 inst_cell_119_86 ( BL86, BLN86, WL119);
sram_cell_6t_3 inst_cell_119_85 ( BL85, BLN85, WL119);
sram_cell_6t_3 inst_cell_119_84 ( BL84, BLN84, WL119);
sram_cell_6t_3 inst_cell_119_83 ( BL83, BLN83, WL119);
sram_cell_6t_3 inst_cell_119_82 ( BL82, BLN82, WL119);
sram_cell_6t_3 inst_cell_119_81 ( BL81, BLN81, WL119);
sram_cell_6t_3 inst_cell_119_80 ( BL80, BLN80, WL119);
sram_cell_6t_3 inst_cell_119_79 ( BL79, BLN79, WL119);
sram_cell_6t_3 inst_cell_119_78 ( BL78, BLN78, WL119);
sram_cell_6t_3 inst_cell_119_77 ( BL77, BLN77, WL119);
sram_cell_6t_3 inst_cell_119_76 ( BL76, BLN76, WL119);
sram_cell_6t_3 inst_cell_119_75 ( BL75, BLN75, WL119);
sram_cell_6t_3 inst_cell_119_74 ( BL74, BLN74, WL119);
sram_cell_6t_3 inst_cell_119_73 ( BL73, BLN73, WL119);
sram_cell_6t_3 inst_cell_119_72 ( BL72, BLN72, WL119);
sram_cell_6t_3 inst_cell_119_71 ( BL71, BLN71, WL119);
sram_cell_6t_3 inst_cell_119_70 ( BL70, BLN70, WL119);
sram_cell_6t_3 inst_cell_119_69 ( BL69, BLN69, WL119);
sram_cell_6t_3 inst_cell_119_68 ( BL68, BLN68, WL119);
sram_cell_6t_3 inst_cell_119_67 ( BL67, BLN67, WL119);
sram_cell_6t_3 inst_cell_119_66 ( BL66, BLN66, WL119);
sram_cell_6t_3 inst_cell_119_65 ( BL65, BLN65, WL119);
sram_cell_6t_3 inst_cell_119_64 ( BL64, BLN64, WL119);
sram_cell_6t_3 inst_cell_119_63 ( BL63, BLN63, WL119);
sram_cell_6t_3 inst_cell_119_62 ( BL62, BLN62, WL119);
sram_cell_6t_3 inst_cell_119_61 ( BL61, BLN61, WL119);
sram_cell_6t_3 inst_cell_119_60 ( BL60, BLN60, WL119);
sram_cell_6t_3 inst_cell_119_59 ( BL59, BLN59, WL119);
sram_cell_6t_3 inst_cell_119_58 ( BL58, BLN58, WL119);
sram_cell_6t_3 inst_cell_119_57 ( BL57, BLN57, WL119);
sram_cell_6t_3 inst_cell_119_56 ( BL56, BLN56, WL119);
sram_cell_6t_3 inst_cell_119_55 ( BL55, BLN55, WL119);
sram_cell_6t_3 inst_cell_119_54 ( BL54, BLN54, WL119);
sram_cell_6t_3 inst_cell_119_53 ( BL53, BLN53, WL119);
sram_cell_6t_3 inst_cell_119_52 ( BL52, BLN52, WL119);
sram_cell_6t_3 inst_cell_119_51 ( BL51, BLN51, WL119);
sram_cell_6t_3 inst_cell_119_50 ( BL50, BLN50, WL119);
sram_cell_6t_3 inst_cell_119_49 ( BL49, BLN49, WL119);
sram_cell_6t_3 inst_cell_119_48 ( BL48, BLN48, WL119);
sram_cell_6t_3 inst_cell_119_47 ( BL47, BLN47, WL119);
sram_cell_6t_3 inst_cell_119_46 ( BL46, BLN46, WL119);
sram_cell_6t_3 inst_cell_119_45 ( BL45, BLN45, WL119);
sram_cell_6t_3 inst_cell_119_44 ( BL44, BLN44, WL119);
sram_cell_6t_3 inst_cell_119_43 ( BL43, BLN43, WL119);
sram_cell_6t_3 inst_cell_119_42 ( BL42, BLN42, WL119);
sram_cell_6t_3 inst_cell_119_41 ( BL41, BLN41, WL119);
sram_cell_6t_3 inst_cell_119_40 ( BL40, BLN40, WL119);
sram_cell_6t_3 inst_cell_119_39 ( BL39, BLN39, WL119);
sram_cell_6t_3 inst_cell_119_38 ( BL38, BLN38, WL119);
sram_cell_6t_3 inst_cell_119_37 ( BL37, BLN37, WL119);
sram_cell_6t_3 inst_cell_119_36 ( BL36, BLN36, WL119);
sram_cell_6t_3 inst_cell_119_35 ( BL35, BLN35, WL119);
sram_cell_6t_3 inst_cell_119_34 ( BL34, BLN34, WL119);
sram_cell_6t_3 inst_cell_119_33 ( BL33, BLN33, WL119);
sram_cell_6t_3 inst_cell_119_32 ( BL32, BLN32, WL119);
sram_cell_6t_3 inst_cell_119_31 ( BL31, BLN31, WL119);
sram_cell_6t_3 inst_cell_119_30 ( BL30, BLN30, WL119);
sram_cell_6t_3 inst_cell_119_29 ( BL29, BLN29, WL119);
sram_cell_6t_3 inst_cell_119_28 ( BL28, BLN28, WL119);
sram_cell_6t_3 inst_cell_119_27 ( BL27, BLN27, WL119);
sram_cell_6t_3 inst_cell_119_26 ( BL26, BLN26, WL119);
sram_cell_6t_3 inst_cell_119_25 ( BL25, BLN25, WL119);
sram_cell_6t_3 inst_cell_119_24 ( BL24, BLN24, WL119);
sram_cell_6t_3 inst_cell_119_23 ( BL23, BLN23, WL119);
sram_cell_6t_3 inst_cell_119_22 ( BL22, BLN22, WL119);
sram_cell_6t_3 inst_cell_119_21 ( BL21, BLN21, WL119);
sram_cell_6t_3 inst_cell_119_20 ( BL20, BLN20, WL119);
sram_cell_6t_3 inst_cell_119_19 ( BL19, BLN19, WL119);
sram_cell_6t_3 inst_cell_119_18 ( BL18, BLN18, WL119);
sram_cell_6t_3 inst_cell_119_17 ( BL17, BLN17, WL119);
sram_cell_6t_3 inst_cell_119_16 ( BL16, BLN16, WL119);
sram_cell_6t_3 inst_cell_119_15 ( BL15, BLN15, WL119);
sram_cell_6t_3 inst_cell_119_14 ( BL14, BLN14, WL119);
sram_cell_6t_3 inst_cell_119_13 ( BL13, BLN13, WL119);
sram_cell_6t_3 inst_cell_119_12 ( BL12, BLN12, WL119);
sram_cell_6t_3 inst_cell_119_11 ( BL11, BLN11, WL119);
sram_cell_6t_3 inst_cell_119_10 ( BL10, BLN10, WL119);
sram_cell_6t_3 inst_cell_119_9 ( BL9, BLN9, WL119);
sram_cell_6t_3 inst_cell_119_8 ( BL8, BLN8, WL119);
sram_cell_6t_3 inst_cell_119_7 ( BL7, BLN7, WL119);
sram_cell_6t_3 inst_cell_119_6 ( BL6, BLN6, WL119);
sram_cell_6t_3 inst_cell_119_5 ( BL5, BLN5, WL119);
sram_cell_6t_3 inst_cell_119_4 ( BL4, BLN4, WL119);
sram_cell_6t_3 inst_cell_119_3 ( BL3, BLN3, WL119);
sram_cell_6t_3 inst_cell_119_2 ( BL2, BLN2, WL119);
sram_cell_6t_3 inst_cell_119_1 ( BL1, BLN1, WL119);
sram_cell_6t_3 inst_cell_119_0 ( BL0, BLN0, WL119);
sram_cell_6t_3 inst_cell_118_127 ( BL127, BLN127, WL118);
sram_cell_6t_3 inst_cell_118_126 ( BL126, BLN126, WL118);
sram_cell_6t_3 inst_cell_118_125 ( BL125, BLN125, WL118);
sram_cell_6t_3 inst_cell_118_124 ( BL124, BLN124, WL118);
sram_cell_6t_3 inst_cell_118_123 ( BL123, BLN123, WL118);
sram_cell_6t_3 inst_cell_118_122 ( BL122, BLN122, WL118);
sram_cell_6t_3 inst_cell_118_121 ( BL121, BLN121, WL118);
sram_cell_6t_3 inst_cell_118_120 ( BL120, BLN120, WL118);
sram_cell_6t_3 inst_cell_118_119 ( BL119, BLN119, WL118);
sram_cell_6t_3 inst_cell_118_118 ( BL118, BLN118, WL118);
sram_cell_6t_3 inst_cell_118_117 ( BL117, BLN117, WL118);
sram_cell_6t_3 inst_cell_118_116 ( BL116, BLN116, WL118);
sram_cell_6t_3 inst_cell_118_115 ( BL115, BLN115, WL118);
sram_cell_6t_3 inst_cell_118_114 ( BL114, BLN114, WL118);
sram_cell_6t_3 inst_cell_118_113 ( BL113, BLN113, WL118);
sram_cell_6t_3 inst_cell_118_112 ( BL112, BLN112, WL118);
sram_cell_6t_3 inst_cell_118_111 ( BL111, BLN111, WL118);
sram_cell_6t_3 inst_cell_118_110 ( BL110, BLN110, WL118);
sram_cell_6t_3 inst_cell_118_109 ( BL109, BLN109, WL118);
sram_cell_6t_3 inst_cell_118_108 ( BL108, BLN108, WL118);
sram_cell_6t_3 inst_cell_118_107 ( BL107, BLN107, WL118);
sram_cell_6t_3 inst_cell_118_106 ( BL106, BLN106, WL118);
sram_cell_6t_3 inst_cell_118_105 ( BL105, BLN105, WL118);
sram_cell_6t_3 inst_cell_118_104 ( BL104, BLN104, WL118);
sram_cell_6t_3 inst_cell_118_103 ( BL103, BLN103, WL118);
sram_cell_6t_3 inst_cell_118_102 ( BL102, BLN102, WL118);
sram_cell_6t_3 inst_cell_118_101 ( BL101, BLN101, WL118);
sram_cell_6t_3 inst_cell_118_100 ( BL100, BLN100, WL118);
sram_cell_6t_3 inst_cell_118_99 ( BL99, BLN99, WL118);
sram_cell_6t_3 inst_cell_118_98 ( BL98, BLN98, WL118);
sram_cell_6t_3 inst_cell_118_97 ( BL97, BLN97, WL118);
sram_cell_6t_3 inst_cell_118_96 ( BL96, BLN96, WL118);
sram_cell_6t_3 inst_cell_118_95 ( BL95, BLN95, WL118);
sram_cell_6t_3 inst_cell_118_94 ( BL94, BLN94, WL118);
sram_cell_6t_3 inst_cell_118_93 ( BL93, BLN93, WL118);
sram_cell_6t_3 inst_cell_118_92 ( BL92, BLN92, WL118);
sram_cell_6t_3 inst_cell_118_91 ( BL91, BLN91, WL118);
sram_cell_6t_3 inst_cell_118_90 ( BL90, BLN90, WL118);
sram_cell_6t_3 inst_cell_118_89 ( BL89, BLN89, WL118);
sram_cell_6t_3 inst_cell_118_88 ( BL88, BLN88, WL118);
sram_cell_6t_3 inst_cell_118_87 ( BL87, BLN87, WL118);
sram_cell_6t_3 inst_cell_118_86 ( BL86, BLN86, WL118);
sram_cell_6t_3 inst_cell_118_85 ( BL85, BLN85, WL118);
sram_cell_6t_3 inst_cell_118_84 ( BL84, BLN84, WL118);
sram_cell_6t_3 inst_cell_118_83 ( BL83, BLN83, WL118);
sram_cell_6t_3 inst_cell_118_82 ( BL82, BLN82, WL118);
sram_cell_6t_3 inst_cell_118_81 ( BL81, BLN81, WL118);
sram_cell_6t_3 inst_cell_118_80 ( BL80, BLN80, WL118);
sram_cell_6t_3 inst_cell_118_79 ( BL79, BLN79, WL118);
sram_cell_6t_3 inst_cell_118_78 ( BL78, BLN78, WL118);
sram_cell_6t_3 inst_cell_118_77 ( BL77, BLN77, WL118);
sram_cell_6t_3 inst_cell_118_76 ( BL76, BLN76, WL118);
sram_cell_6t_3 inst_cell_118_75 ( BL75, BLN75, WL118);
sram_cell_6t_3 inst_cell_118_74 ( BL74, BLN74, WL118);
sram_cell_6t_3 inst_cell_118_73 ( BL73, BLN73, WL118);
sram_cell_6t_3 inst_cell_118_72 ( BL72, BLN72, WL118);
sram_cell_6t_3 inst_cell_118_71 ( BL71, BLN71, WL118);
sram_cell_6t_3 inst_cell_118_70 ( BL70, BLN70, WL118);
sram_cell_6t_3 inst_cell_118_69 ( BL69, BLN69, WL118);
sram_cell_6t_3 inst_cell_118_68 ( BL68, BLN68, WL118);
sram_cell_6t_3 inst_cell_118_67 ( BL67, BLN67, WL118);
sram_cell_6t_3 inst_cell_118_66 ( BL66, BLN66, WL118);
sram_cell_6t_3 inst_cell_118_65 ( BL65, BLN65, WL118);
sram_cell_6t_3 inst_cell_118_64 ( BL64, BLN64, WL118);
sram_cell_6t_3 inst_cell_118_63 ( BL63, BLN63, WL118);
sram_cell_6t_3 inst_cell_118_62 ( BL62, BLN62, WL118);
sram_cell_6t_3 inst_cell_118_61 ( BL61, BLN61, WL118);
sram_cell_6t_3 inst_cell_118_60 ( BL60, BLN60, WL118);
sram_cell_6t_3 inst_cell_118_59 ( BL59, BLN59, WL118);
sram_cell_6t_3 inst_cell_118_58 ( BL58, BLN58, WL118);
sram_cell_6t_3 inst_cell_118_57 ( BL57, BLN57, WL118);
sram_cell_6t_3 inst_cell_118_56 ( BL56, BLN56, WL118);
sram_cell_6t_3 inst_cell_118_55 ( BL55, BLN55, WL118);
sram_cell_6t_3 inst_cell_118_54 ( BL54, BLN54, WL118);
sram_cell_6t_3 inst_cell_118_53 ( BL53, BLN53, WL118);
sram_cell_6t_3 inst_cell_118_52 ( BL52, BLN52, WL118);
sram_cell_6t_3 inst_cell_118_51 ( BL51, BLN51, WL118);
sram_cell_6t_3 inst_cell_118_50 ( BL50, BLN50, WL118);
sram_cell_6t_3 inst_cell_118_49 ( BL49, BLN49, WL118);
sram_cell_6t_3 inst_cell_118_48 ( BL48, BLN48, WL118);
sram_cell_6t_3 inst_cell_118_47 ( BL47, BLN47, WL118);
sram_cell_6t_3 inst_cell_118_46 ( BL46, BLN46, WL118);
sram_cell_6t_3 inst_cell_118_45 ( BL45, BLN45, WL118);
sram_cell_6t_3 inst_cell_118_44 ( BL44, BLN44, WL118);
sram_cell_6t_3 inst_cell_118_43 ( BL43, BLN43, WL118);
sram_cell_6t_3 inst_cell_118_42 ( BL42, BLN42, WL118);
sram_cell_6t_3 inst_cell_118_41 ( BL41, BLN41, WL118);
sram_cell_6t_3 inst_cell_118_40 ( BL40, BLN40, WL118);
sram_cell_6t_3 inst_cell_118_39 ( BL39, BLN39, WL118);
sram_cell_6t_3 inst_cell_118_38 ( BL38, BLN38, WL118);
sram_cell_6t_3 inst_cell_118_37 ( BL37, BLN37, WL118);
sram_cell_6t_3 inst_cell_118_36 ( BL36, BLN36, WL118);
sram_cell_6t_3 inst_cell_118_35 ( BL35, BLN35, WL118);
sram_cell_6t_3 inst_cell_118_34 ( BL34, BLN34, WL118);
sram_cell_6t_3 inst_cell_118_33 ( BL33, BLN33, WL118);
sram_cell_6t_3 inst_cell_118_32 ( BL32, BLN32, WL118);
sram_cell_6t_3 inst_cell_118_31 ( BL31, BLN31, WL118);
sram_cell_6t_3 inst_cell_118_30 ( BL30, BLN30, WL118);
sram_cell_6t_3 inst_cell_118_29 ( BL29, BLN29, WL118);
sram_cell_6t_3 inst_cell_118_28 ( BL28, BLN28, WL118);
sram_cell_6t_3 inst_cell_118_27 ( BL27, BLN27, WL118);
sram_cell_6t_3 inst_cell_118_26 ( BL26, BLN26, WL118);
sram_cell_6t_3 inst_cell_118_25 ( BL25, BLN25, WL118);
sram_cell_6t_3 inst_cell_118_24 ( BL24, BLN24, WL118);
sram_cell_6t_3 inst_cell_118_23 ( BL23, BLN23, WL118);
sram_cell_6t_3 inst_cell_118_22 ( BL22, BLN22, WL118);
sram_cell_6t_3 inst_cell_118_21 ( BL21, BLN21, WL118);
sram_cell_6t_3 inst_cell_118_20 ( BL20, BLN20, WL118);
sram_cell_6t_3 inst_cell_118_19 ( BL19, BLN19, WL118);
sram_cell_6t_3 inst_cell_118_18 ( BL18, BLN18, WL118);
sram_cell_6t_3 inst_cell_118_17 ( BL17, BLN17, WL118);
sram_cell_6t_3 inst_cell_118_16 ( BL16, BLN16, WL118);
sram_cell_6t_3 inst_cell_118_15 ( BL15, BLN15, WL118);
sram_cell_6t_3 inst_cell_118_14 ( BL14, BLN14, WL118);
sram_cell_6t_3 inst_cell_118_13 ( BL13, BLN13, WL118);
sram_cell_6t_3 inst_cell_118_12 ( BL12, BLN12, WL118);
sram_cell_6t_3 inst_cell_118_11 ( BL11, BLN11, WL118);
sram_cell_6t_3 inst_cell_118_10 ( BL10, BLN10, WL118);
sram_cell_6t_3 inst_cell_118_9 ( BL9, BLN9, WL118);
sram_cell_6t_3 inst_cell_118_8 ( BL8, BLN8, WL118);
sram_cell_6t_3 inst_cell_118_7 ( BL7, BLN7, WL118);
sram_cell_6t_3 inst_cell_118_6 ( BL6, BLN6, WL118);
sram_cell_6t_3 inst_cell_118_5 ( BL5, BLN5, WL118);
sram_cell_6t_3 inst_cell_118_4 ( BL4, BLN4, WL118);
sram_cell_6t_3 inst_cell_118_3 ( BL3, BLN3, WL118);
sram_cell_6t_3 inst_cell_118_2 ( BL2, BLN2, WL118);
sram_cell_6t_3 inst_cell_118_1 ( BL1, BLN1, WL118);
sram_cell_6t_3 inst_cell_118_0 ( BL0, BLN0, WL118);
sram_cell_6t_3 inst_cell_117_127 ( BL127, BLN127, WL117);
sram_cell_6t_3 inst_cell_117_126 ( BL126, BLN126, WL117);
sram_cell_6t_3 inst_cell_117_125 ( BL125, BLN125, WL117);
sram_cell_6t_3 inst_cell_117_124 ( BL124, BLN124, WL117);
sram_cell_6t_3 inst_cell_117_123 ( BL123, BLN123, WL117);
sram_cell_6t_3 inst_cell_117_122 ( BL122, BLN122, WL117);
sram_cell_6t_3 inst_cell_117_121 ( BL121, BLN121, WL117);
sram_cell_6t_3 inst_cell_117_120 ( BL120, BLN120, WL117);
sram_cell_6t_3 inst_cell_117_119 ( BL119, BLN119, WL117);
sram_cell_6t_3 inst_cell_117_118 ( BL118, BLN118, WL117);
sram_cell_6t_3 inst_cell_117_117 ( BL117, BLN117, WL117);
sram_cell_6t_3 inst_cell_117_116 ( BL116, BLN116, WL117);
sram_cell_6t_3 inst_cell_117_115 ( BL115, BLN115, WL117);
sram_cell_6t_3 inst_cell_117_114 ( BL114, BLN114, WL117);
sram_cell_6t_3 inst_cell_117_113 ( BL113, BLN113, WL117);
sram_cell_6t_3 inst_cell_117_112 ( BL112, BLN112, WL117);
sram_cell_6t_3 inst_cell_117_111 ( BL111, BLN111, WL117);
sram_cell_6t_3 inst_cell_117_110 ( BL110, BLN110, WL117);
sram_cell_6t_3 inst_cell_117_109 ( BL109, BLN109, WL117);
sram_cell_6t_3 inst_cell_117_108 ( BL108, BLN108, WL117);
sram_cell_6t_3 inst_cell_117_107 ( BL107, BLN107, WL117);
sram_cell_6t_3 inst_cell_117_106 ( BL106, BLN106, WL117);
sram_cell_6t_3 inst_cell_117_105 ( BL105, BLN105, WL117);
sram_cell_6t_3 inst_cell_117_104 ( BL104, BLN104, WL117);
sram_cell_6t_3 inst_cell_117_103 ( BL103, BLN103, WL117);
sram_cell_6t_3 inst_cell_117_102 ( BL102, BLN102, WL117);
sram_cell_6t_3 inst_cell_117_101 ( BL101, BLN101, WL117);
sram_cell_6t_3 inst_cell_117_100 ( BL100, BLN100, WL117);
sram_cell_6t_3 inst_cell_117_99 ( BL99, BLN99, WL117);
sram_cell_6t_3 inst_cell_117_98 ( BL98, BLN98, WL117);
sram_cell_6t_3 inst_cell_117_97 ( BL97, BLN97, WL117);
sram_cell_6t_3 inst_cell_117_96 ( BL96, BLN96, WL117);
sram_cell_6t_3 inst_cell_117_95 ( BL95, BLN95, WL117);
sram_cell_6t_3 inst_cell_117_94 ( BL94, BLN94, WL117);
sram_cell_6t_3 inst_cell_117_93 ( BL93, BLN93, WL117);
sram_cell_6t_3 inst_cell_117_92 ( BL92, BLN92, WL117);
sram_cell_6t_3 inst_cell_117_91 ( BL91, BLN91, WL117);
sram_cell_6t_3 inst_cell_117_90 ( BL90, BLN90, WL117);
sram_cell_6t_3 inst_cell_117_89 ( BL89, BLN89, WL117);
sram_cell_6t_3 inst_cell_117_88 ( BL88, BLN88, WL117);
sram_cell_6t_3 inst_cell_117_87 ( BL87, BLN87, WL117);
sram_cell_6t_3 inst_cell_117_86 ( BL86, BLN86, WL117);
sram_cell_6t_3 inst_cell_117_85 ( BL85, BLN85, WL117);
sram_cell_6t_3 inst_cell_117_84 ( BL84, BLN84, WL117);
sram_cell_6t_3 inst_cell_117_83 ( BL83, BLN83, WL117);
sram_cell_6t_3 inst_cell_117_82 ( BL82, BLN82, WL117);
sram_cell_6t_3 inst_cell_117_81 ( BL81, BLN81, WL117);
sram_cell_6t_3 inst_cell_117_80 ( BL80, BLN80, WL117);
sram_cell_6t_3 inst_cell_117_79 ( BL79, BLN79, WL117);
sram_cell_6t_3 inst_cell_117_78 ( BL78, BLN78, WL117);
sram_cell_6t_3 inst_cell_117_77 ( BL77, BLN77, WL117);
sram_cell_6t_3 inst_cell_117_76 ( BL76, BLN76, WL117);
sram_cell_6t_3 inst_cell_117_75 ( BL75, BLN75, WL117);
sram_cell_6t_3 inst_cell_117_74 ( BL74, BLN74, WL117);
sram_cell_6t_3 inst_cell_117_73 ( BL73, BLN73, WL117);
sram_cell_6t_3 inst_cell_117_72 ( BL72, BLN72, WL117);
sram_cell_6t_3 inst_cell_117_71 ( BL71, BLN71, WL117);
sram_cell_6t_3 inst_cell_117_70 ( BL70, BLN70, WL117);
sram_cell_6t_3 inst_cell_117_69 ( BL69, BLN69, WL117);
sram_cell_6t_3 inst_cell_117_68 ( BL68, BLN68, WL117);
sram_cell_6t_3 inst_cell_117_67 ( BL67, BLN67, WL117);
sram_cell_6t_3 inst_cell_117_66 ( BL66, BLN66, WL117);
sram_cell_6t_3 inst_cell_117_65 ( BL65, BLN65, WL117);
sram_cell_6t_3 inst_cell_117_64 ( BL64, BLN64, WL117);
sram_cell_6t_3 inst_cell_117_63 ( BL63, BLN63, WL117);
sram_cell_6t_3 inst_cell_117_62 ( BL62, BLN62, WL117);
sram_cell_6t_3 inst_cell_117_61 ( BL61, BLN61, WL117);
sram_cell_6t_3 inst_cell_117_60 ( BL60, BLN60, WL117);
sram_cell_6t_3 inst_cell_117_59 ( BL59, BLN59, WL117);
sram_cell_6t_3 inst_cell_117_58 ( BL58, BLN58, WL117);
sram_cell_6t_3 inst_cell_117_57 ( BL57, BLN57, WL117);
sram_cell_6t_3 inst_cell_117_56 ( BL56, BLN56, WL117);
sram_cell_6t_3 inst_cell_117_55 ( BL55, BLN55, WL117);
sram_cell_6t_3 inst_cell_117_54 ( BL54, BLN54, WL117);
sram_cell_6t_3 inst_cell_117_53 ( BL53, BLN53, WL117);
sram_cell_6t_3 inst_cell_117_52 ( BL52, BLN52, WL117);
sram_cell_6t_3 inst_cell_117_51 ( BL51, BLN51, WL117);
sram_cell_6t_3 inst_cell_117_50 ( BL50, BLN50, WL117);
sram_cell_6t_3 inst_cell_117_49 ( BL49, BLN49, WL117);
sram_cell_6t_3 inst_cell_117_48 ( BL48, BLN48, WL117);
sram_cell_6t_3 inst_cell_117_47 ( BL47, BLN47, WL117);
sram_cell_6t_3 inst_cell_117_46 ( BL46, BLN46, WL117);
sram_cell_6t_3 inst_cell_117_45 ( BL45, BLN45, WL117);
sram_cell_6t_3 inst_cell_117_44 ( BL44, BLN44, WL117);
sram_cell_6t_3 inst_cell_117_43 ( BL43, BLN43, WL117);
sram_cell_6t_3 inst_cell_117_42 ( BL42, BLN42, WL117);
sram_cell_6t_3 inst_cell_117_41 ( BL41, BLN41, WL117);
sram_cell_6t_3 inst_cell_117_40 ( BL40, BLN40, WL117);
sram_cell_6t_3 inst_cell_117_39 ( BL39, BLN39, WL117);
sram_cell_6t_3 inst_cell_117_38 ( BL38, BLN38, WL117);
sram_cell_6t_3 inst_cell_117_37 ( BL37, BLN37, WL117);
sram_cell_6t_3 inst_cell_117_36 ( BL36, BLN36, WL117);
sram_cell_6t_3 inst_cell_117_35 ( BL35, BLN35, WL117);
sram_cell_6t_3 inst_cell_117_34 ( BL34, BLN34, WL117);
sram_cell_6t_3 inst_cell_117_33 ( BL33, BLN33, WL117);
sram_cell_6t_3 inst_cell_117_32 ( BL32, BLN32, WL117);
sram_cell_6t_3 inst_cell_117_31 ( BL31, BLN31, WL117);
sram_cell_6t_3 inst_cell_117_30 ( BL30, BLN30, WL117);
sram_cell_6t_3 inst_cell_117_29 ( BL29, BLN29, WL117);
sram_cell_6t_3 inst_cell_117_28 ( BL28, BLN28, WL117);
sram_cell_6t_3 inst_cell_117_27 ( BL27, BLN27, WL117);
sram_cell_6t_3 inst_cell_117_26 ( BL26, BLN26, WL117);
sram_cell_6t_3 inst_cell_117_25 ( BL25, BLN25, WL117);
sram_cell_6t_3 inst_cell_117_24 ( BL24, BLN24, WL117);
sram_cell_6t_3 inst_cell_117_23 ( BL23, BLN23, WL117);
sram_cell_6t_3 inst_cell_117_22 ( BL22, BLN22, WL117);
sram_cell_6t_3 inst_cell_117_21 ( BL21, BLN21, WL117);
sram_cell_6t_3 inst_cell_117_20 ( BL20, BLN20, WL117);
sram_cell_6t_3 inst_cell_117_19 ( BL19, BLN19, WL117);
sram_cell_6t_3 inst_cell_117_18 ( BL18, BLN18, WL117);
sram_cell_6t_3 inst_cell_117_17 ( BL17, BLN17, WL117);
sram_cell_6t_3 inst_cell_117_16 ( BL16, BLN16, WL117);
sram_cell_6t_3 inst_cell_117_15 ( BL15, BLN15, WL117);
sram_cell_6t_3 inst_cell_117_14 ( BL14, BLN14, WL117);
sram_cell_6t_3 inst_cell_117_13 ( BL13, BLN13, WL117);
sram_cell_6t_3 inst_cell_117_12 ( BL12, BLN12, WL117);
sram_cell_6t_3 inst_cell_117_11 ( BL11, BLN11, WL117);
sram_cell_6t_3 inst_cell_117_10 ( BL10, BLN10, WL117);
sram_cell_6t_3 inst_cell_117_9 ( BL9, BLN9, WL117);
sram_cell_6t_3 inst_cell_117_8 ( BL8, BLN8, WL117);
sram_cell_6t_3 inst_cell_117_7 ( BL7, BLN7, WL117);
sram_cell_6t_3 inst_cell_117_6 ( BL6, BLN6, WL117);
sram_cell_6t_3 inst_cell_117_5 ( BL5, BLN5, WL117);
sram_cell_6t_3 inst_cell_117_4 ( BL4, BLN4, WL117);
sram_cell_6t_3 inst_cell_117_3 ( BL3, BLN3, WL117);
sram_cell_6t_3 inst_cell_117_2 ( BL2, BLN2, WL117);
sram_cell_6t_3 inst_cell_117_1 ( BL1, BLN1, WL117);
sram_cell_6t_3 inst_cell_117_0 ( BL0, BLN0, WL117);
sram_cell_6t_3 inst_cell_116_127 ( BL127, BLN127, WL116);
sram_cell_6t_3 inst_cell_116_126 ( BL126, BLN126, WL116);
sram_cell_6t_3 inst_cell_116_125 ( BL125, BLN125, WL116);
sram_cell_6t_3 inst_cell_116_124 ( BL124, BLN124, WL116);
sram_cell_6t_3 inst_cell_116_123 ( BL123, BLN123, WL116);
sram_cell_6t_3 inst_cell_116_122 ( BL122, BLN122, WL116);
sram_cell_6t_3 inst_cell_116_121 ( BL121, BLN121, WL116);
sram_cell_6t_3 inst_cell_116_120 ( BL120, BLN120, WL116);
sram_cell_6t_3 inst_cell_116_119 ( BL119, BLN119, WL116);
sram_cell_6t_3 inst_cell_116_118 ( BL118, BLN118, WL116);
sram_cell_6t_3 inst_cell_116_117 ( BL117, BLN117, WL116);
sram_cell_6t_3 inst_cell_116_116 ( BL116, BLN116, WL116);
sram_cell_6t_3 inst_cell_116_115 ( BL115, BLN115, WL116);
sram_cell_6t_3 inst_cell_116_114 ( BL114, BLN114, WL116);
sram_cell_6t_3 inst_cell_116_113 ( BL113, BLN113, WL116);
sram_cell_6t_3 inst_cell_116_112 ( BL112, BLN112, WL116);
sram_cell_6t_3 inst_cell_116_111 ( BL111, BLN111, WL116);
sram_cell_6t_3 inst_cell_116_110 ( BL110, BLN110, WL116);
sram_cell_6t_3 inst_cell_116_109 ( BL109, BLN109, WL116);
sram_cell_6t_3 inst_cell_116_108 ( BL108, BLN108, WL116);
sram_cell_6t_3 inst_cell_116_107 ( BL107, BLN107, WL116);
sram_cell_6t_3 inst_cell_116_106 ( BL106, BLN106, WL116);
sram_cell_6t_3 inst_cell_116_105 ( BL105, BLN105, WL116);
sram_cell_6t_3 inst_cell_116_104 ( BL104, BLN104, WL116);
sram_cell_6t_3 inst_cell_116_103 ( BL103, BLN103, WL116);
sram_cell_6t_3 inst_cell_116_102 ( BL102, BLN102, WL116);
sram_cell_6t_3 inst_cell_116_101 ( BL101, BLN101, WL116);
sram_cell_6t_3 inst_cell_116_100 ( BL100, BLN100, WL116);
sram_cell_6t_3 inst_cell_116_99 ( BL99, BLN99, WL116);
sram_cell_6t_3 inst_cell_116_98 ( BL98, BLN98, WL116);
sram_cell_6t_3 inst_cell_116_97 ( BL97, BLN97, WL116);
sram_cell_6t_3 inst_cell_116_96 ( BL96, BLN96, WL116);
sram_cell_6t_3 inst_cell_116_95 ( BL95, BLN95, WL116);
sram_cell_6t_3 inst_cell_116_94 ( BL94, BLN94, WL116);
sram_cell_6t_3 inst_cell_116_93 ( BL93, BLN93, WL116);
sram_cell_6t_3 inst_cell_116_92 ( BL92, BLN92, WL116);
sram_cell_6t_3 inst_cell_116_91 ( BL91, BLN91, WL116);
sram_cell_6t_3 inst_cell_116_90 ( BL90, BLN90, WL116);
sram_cell_6t_3 inst_cell_116_89 ( BL89, BLN89, WL116);
sram_cell_6t_3 inst_cell_116_88 ( BL88, BLN88, WL116);
sram_cell_6t_3 inst_cell_116_87 ( BL87, BLN87, WL116);
sram_cell_6t_3 inst_cell_116_86 ( BL86, BLN86, WL116);
sram_cell_6t_3 inst_cell_116_85 ( BL85, BLN85, WL116);
sram_cell_6t_3 inst_cell_116_84 ( BL84, BLN84, WL116);
sram_cell_6t_3 inst_cell_116_83 ( BL83, BLN83, WL116);
sram_cell_6t_3 inst_cell_116_82 ( BL82, BLN82, WL116);
sram_cell_6t_3 inst_cell_116_81 ( BL81, BLN81, WL116);
sram_cell_6t_3 inst_cell_116_80 ( BL80, BLN80, WL116);
sram_cell_6t_3 inst_cell_116_79 ( BL79, BLN79, WL116);
sram_cell_6t_3 inst_cell_116_78 ( BL78, BLN78, WL116);
sram_cell_6t_3 inst_cell_116_77 ( BL77, BLN77, WL116);
sram_cell_6t_3 inst_cell_116_76 ( BL76, BLN76, WL116);
sram_cell_6t_3 inst_cell_116_75 ( BL75, BLN75, WL116);
sram_cell_6t_3 inst_cell_116_74 ( BL74, BLN74, WL116);
sram_cell_6t_3 inst_cell_116_73 ( BL73, BLN73, WL116);
sram_cell_6t_3 inst_cell_116_72 ( BL72, BLN72, WL116);
sram_cell_6t_3 inst_cell_116_71 ( BL71, BLN71, WL116);
sram_cell_6t_3 inst_cell_116_70 ( BL70, BLN70, WL116);
sram_cell_6t_3 inst_cell_116_69 ( BL69, BLN69, WL116);
sram_cell_6t_3 inst_cell_116_68 ( BL68, BLN68, WL116);
sram_cell_6t_3 inst_cell_116_67 ( BL67, BLN67, WL116);
sram_cell_6t_3 inst_cell_116_66 ( BL66, BLN66, WL116);
sram_cell_6t_3 inst_cell_116_65 ( BL65, BLN65, WL116);
sram_cell_6t_3 inst_cell_116_64 ( BL64, BLN64, WL116);
sram_cell_6t_3 inst_cell_116_63 ( BL63, BLN63, WL116);
sram_cell_6t_3 inst_cell_116_62 ( BL62, BLN62, WL116);
sram_cell_6t_3 inst_cell_116_61 ( BL61, BLN61, WL116);
sram_cell_6t_3 inst_cell_116_60 ( BL60, BLN60, WL116);
sram_cell_6t_3 inst_cell_116_59 ( BL59, BLN59, WL116);
sram_cell_6t_3 inst_cell_116_58 ( BL58, BLN58, WL116);
sram_cell_6t_3 inst_cell_116_57 ( BL57, BLN57, WL116);
sram_cell_6t_3 inst_cell_116_56 ( BL56, BLN56, WL116);
sram_cell_6t_3 inst_cell_116_55 ( BL55, BLN55, WL116);
sram_cell_6t_3 inst_cell_116_54 ( BL54, BLN54, WL116);
sram_cell_6t_3 inst_cell_116_53 ( BL53, BLN53, WL116);
sram_cell_6t_3 inst_cell_116_52 ( BL52, BLN52, WL116);
sram_cell_6t_3 inst_cell_116_51 ( BL51, BLN51, WL116);
sram_cell_6t_3 inst_cell_116_50 ( BL50, BLN50, WL116);
sram_cell_6t_3 inst_cell_116_49 ( BL49, BLN49, WL116);
sram_cell_6t_3 inst_cell_116_48 ( BL48, BLN48, WL116);
sram_cell_6t_3 inst_cell_116_47 ( BL47, BLN47, WL116);
sram_cell_6t_3 inst_cell_116_46 ( BL46, BLN46, WL116);
sram_cell_6t_3 inst_cell_116_45 ( BL45, BLN45, WL116);
sram_cell_6t_3 inst_cell_116_44 ( BL44, BLN44, WL116);
sram_cell_6t_3 inst_cell_116_43 ( BL43, BLN43, WL116);
sram_cell_6t_3 inst_cell_116_42 ( BL42, BLN42, WL116);
sram_cell_6t_3 inst_cell_116_41 ( BL41, BLN41, WL116);
sram_cell_6t_3 inst_cell_116_40 ( BL40, BLN40, WL116);
sram_cell_6t_3 inst_cell_116_39 ( BL39, BLN39, WL116);
sram_cell_6t_3 inst_cell_116_38 ( BL38, BLN38, WL116);
sram_cell_6t_3 inst_cell_116_37 ( BL37, BLN37, WL116);
sram_cell_6t_3 inst_cell_116_36 ( BL36, BLN36, WL116);
sram_cell_6t_3 inst_cell_116_35 ( BL35, BLN35, WL116);
sram_cell_6t_3 inst_cell_116_34 ( BL34, BLN34, WL116);
sram_cell_6t_3 inst_cell_116_33 ( BL33, BLN33, WL116);
sram_cell_6t_3 inst_cell_116_32 ( BL32, BLN32, WL116);
sram_cell_6t_3 inst_cell_116_31 ( BL31, BLN31, WL116);
sram_cell_6t_3 inst_cell_116_30 ( BL30, BLN30, WL116);
sram_cell_6t_3 inst_cell_116_29 ( BL29, BLN29, WL116);
sram_cell_6t_3 inst_cell_116_28 ( BL28, BLN28, WL116);
sram_cell_6t_3 inst_cell_116_27 ( BL27, BLN27, WL116);
sram_cell_6t_3 inst_cell_116_26 ( BL26, BLN26, WL116);
sram_cell_6t_3 inst_cell_116_25 ( BL25, BLN25, WL116);
sram_cell_6t_3 inst_cell_116_24 ( BL24, BLN24, WL116);
sram_cell_6t_3 inst_cell_116_23 ( BL23, BLN23, WL116);
sram_cell_6t_3 inst_cell_116_22 ( BL22, BLN22, WL116);
sram_cell_6t_3 inst_cell_116_21 ( BL21, BLN21, WL116);
sram_cell_6t_3 inst_cell_116_20 ( BL20, BLN20, WL116);
sram_cell_6t_3 inst_cell_116_19 ( BL19, BLN19, WL116);
sram_cell_6t_3 inst_cell_116_18 ( BL18, BLN18, WL116);
sram_cell_6t_3 inst_cell_116_17 ( BL17, BLN17, WL116);
sram_cell_6t_3 inst_cell_116_16 ( BL16, BLN16, WL116);
sram_cell_6t_3 inst_cell_116_15 ( BL15, BLN15, WL116);
sram_cell_6t_3 inst_cell_116_14 ( BL14, BLN14, WL116);
sram_cell_6t_3 inst_cell_116_13 ( BL13, BLN13, WL116);
sram_cell_6t_3 inst_cell_116_12 ( BL12, BLN12, WL116);
sram_cell_6t_3 inst_cell_116_11 ( BL11, BLN11, WL116);
sram_cell_6t_3 inst_cell_116_10 ( BL10, BLN10, WL116);
sram_cell_6t_3 inst_cell_116_9 ( BL9, BLN9, WL116);
sram_cell_6t_3 inst_cell_116_8 ( BL8, BLN8, WL116);
sram_cell_6t_3 inst_cell_116_7 ( BL7, BLN7, WL116);
sram_cell_6t_3 inst_cell_116_6 ( BL6, BLN6, WL116);
sram_cell_6t_3 inst_cell_116_5 ( BL5, BLN5, WL116);
sram_cell_6t_3 inst_cell_116_4 ( BL4, BLN4, WL116);
sram_cell_6t_3 inst_cell_116_3 ( BL3, BLN3, WL116);
sram_cell_6t_3 inst_cell_116_2 ( BL2, BLN2, WL116);
sram_cell_6t_3 inst_cell_116_1 ( BL1, BLN1, WL116);
sram_cell_6t_3 inst_cell_116_0 ( BL0, BLN0, WL116);
sram_cell_6t_3 inst_cell_115_127 ( BL127, BLN127, WL115);
sram_cell_6t_3 inst_cell_115_126 ( BL126, BLN126, WL115);
sram_cell_6t_3 inst_cell_115_125 ( BL125, BLN125, WL115);
sram_cell_6t_3 inst_cell_115_124 ( BL124, BLN124, WL115);
sram_cell_6t_3 inst_cell_115_123 ( BL123, BLN123, WL115);
sram_cell_6t_3 inst_cell_115_122 ( BL122, BLN122, WL115);
sram_cell_6t_3 inst_cell_115_121 ( BL121, BLN121, WL115);
sram_cell_6t_3 inst_cell_115_120 ( BL120, BLN120, WL115);
sram_cell_6t_3 inst_cell_115_119 ( BL119, BLN119, WL115);
sram_cell_6t_3 inst_cell_115_118 ( BL118, BLN118, WL115);
sram_cell_6t_3 inst_cell_115_117 ( BL117, BLN117, WL115);
sram_cell_6t_3 inst_cell_115_116 ( BL116, BLN116, WL115);
sram_cell_6t_3 inst_cell_115_115 ( BL115, BLN115, WL115);
sram_cell_6t_3 inst_cell_115_114 ( BL114, BLN114, WL115);
sram_cell_6t_3 inst_cell_115_113 ( BL113, BLN113, WL115);
sram_cell_6t_3 inst_cell_115_112 ( BL112, BLN112, WL115);
sram_cell_6t_3 inst_cell_115_111 ( BL111, BLN111, WL115);
sram_cell_6t_3 inst_cell_115_110 ( BL110, BLN110, WL115);
sram_cell_6t_3 inst_cell_115_109 ( BL109, BLN109, WL115);
sram_cell_6t_3 inst_cell_115_108 ( BL108, BLN108, WL115);
sram_cell_6t_3 inst_cell_115_107 ( BL107, BLN107, WL115);
sram_cell_6t_3 inst_cell_115_106 ( BL106, BLN106, WL115);
sram_cell_6t_3 inst_cell_115_105 ( BL105, BLN105, WL115);
sram_cell_6t_3 inst_cell_115_104 ( BL104, BLN104, WL115);
sram_cell_6t_3 inst_cell_115_103 ( BL103, BLN103, WL115);
sram_cell_6t_3 inst_cell_115_102 ( BL102, BLN102, WL115);
sram_cell_6t_3 inst_cell_115_101 ( BL101, BLN101, WL115);
sram_cell_6t_3 inst_cell_115_100 ( BL100, BLN100, WL115);
sram_cell_6t_3 inst_cell_115_99 ( BL99, BLN99, WL115);
sram_cell_6t_3 inst_cell_115_98 ( BL98, BLN98, WL115);
sram_cell_6t_3 inst_cell_115_97 ( BL97, BLN97, WL115);
sram_cell_6t_3 inst_cell_115_96 ( BL96, BLN96, WL115);
sram_cell_6t_3 inst_cell_115_95 ( BL95, BLN95, WL115);
sram_cell_6t_3 inst_cell_115_94 ( BL94, BLN94, WL115);
sram_cell_6t_3 inst_cell_115_93 ( BL93, BLN93, WL115);
sram_cell_6t_3 inst_cell_115_92 ( BL92, BLN92, WL115);
sram_cell_6t_3 inst_cell_115_91 ( BL91, BLN91, WL115);
sram_cell_6t_3 inst_cell_115_90 ( BL90, BLN90, WL115);
sram_cell_6t_3 inst_cell_115_89 ( BL89, BLN89, WL115);
sram_cell_6t_3 inst_cell_115_88 ( BL88, BLN88, WL115);
sram_cell_6t_3 inst_cell_115_87 ( BL87, BLN87, WL115);
sram_cell_6t_3 inst_cell_115_86 ( BL86, BLN86, WL115);
sram_cell_6t_3 inst_cell_115_85 ( BL85, BLN85, WL115);
sram_cell_6t_3 inst_cell_115_84 ( BL84, BLN84, WL115);
sram_cell_6t_3 inst_cell_115_83 ( BL83, BLN83, WL115);
sram_cell_6t_3 inst_cell_115_82 ( BL82, BLN82, WL115);
sram_cell_6t_3 inst_cell_115_81 ( BL81, BLN81, WL115);
sram_cell_6t_3 inst_cell_115_80 ( BL80, BLN80, WL115);
sram_cell_6t_3 inst_cell_115_79 ( BL79, BLN79, WL115);
sram_cell_6t_3 inst_cell_115_78 ( BL78, BLN78, WL115);
sram_cell_6t_3 inst_cell_115_77 ( BL77, BLN77, WL115);
sram_cell_6t_3 inst_cell_115_76 ( BL76, BLN76, WL115);
sram_cell_6t_3 inst_cell_115_75 ( BL75, BLN75, WL115);
sram_cell_6t_3 inst_cell_115_74 ( BL74, BLN74, WL115);
sram_cell_6t_3 inst_cell_115_73 ( BL73, BLN73, WL115);
sram_cell_6t_3 inst_cell_115_72 ( BL72, BLN72, WL115);
sram_cell_6t_3 inst_cell_115_71 ( BL71, BLN71, WL115);
sram_cell_6t_3 inst_cell_115_70 ( BL70, BLN70, WL115);
sram_cell_6t_3 inst_cell_115_69 ( BL69, BLN69, WL115);
sram_cell_6t_3 inst_cell_115_68 ( BL68, BLN68, WL115);
sram_cell_6t_3 inst_cell_115_67 ( BL67, BLN67, WL115);
sram_cell_6t_3 inst_cell_115_66 ( BL66, BLN66, WL115);
sram_cell_6t_3 inst_cell_115_65 ( BL65, BLN65, WL115);
sram_cell_6t_3 inst_cell_115_64 ( BL64, BLN64, WL115);
sram_cell_6t_3 inst_cell_115_63 ( BL63, BLN63, WL115);
sram_cell_6t_3 inst_cell_115_62 ( BL62, BLN62, WL115);
sram_cell_6t_3 inst_cell_115_61 ( BL61, BLN61, WL115);
sram_cell_6t_3 inst_cell_115_60 ( BL60, BLN60, WL115);
sram_cell_6t_3 inst_cell_115_59 ( BL59, BLN59, WL115);
sram_cell_6t_3 inst_cell_115_58 ( BL58, BLN58, WL115);
sram_cell_6t_3 inst_cell_115_57 ( BL57, BLN57, WL115);
sram_cell_6t_3 inst_cell_115_56 ( BL56, BLN56, WL115);
sram_cell_6t_3 inst_cell_115_55 ( BL55, BLN55, WL115);
sram_cell_6t_3 inst_cell_115_54 ( BL54, BLN54, WL115);
sram_cell_6t_3 inst_cell_115_53 ( BL53, BLN53, WL115);
sram_cell_6t_3 inst_cell_115_52 ( BL52, BLN52, WL115);
sram_cell_6t_3 inst_cell_115_51 ( BL51, BLN51, WL115);
sram_cell_6t_3 inst_cell_115_50 ( BL50, BLN50, WL115);
sram_cell_6t_3 inst_cell_115_49 ( BL49, BLN49, WL115);
sram_cell_6t_3 inst_cell_115_48 ( BL48, BLN48, WL115);
sram_cell_6t_3 inst_cell_115_47 ( BL47, BLN47, WL115);
sram_cell_6t_3 inst_cell_115_46 ( BL46, BLN46, WL115);
sram_cell_6t_3 inst_cell_115_45 ( BL45, BLN45, WL115);
sram_cell_6t_3 inst_cell_115_44 ( BL44, BLN44, WL115);
sram_cell_6t_3 inst_cell_115_43 ( BL43, BLN43, WL115);
sram_cell_6t_3 inst_cell_115_42 ( BL42, BLN42, WL115);
sram_cell_6t_3 inst_cell_115_41 ( BL41, BLN41, WL115);
sram_cell_6t_3 inst_cell_115_40 ( BL40, BLN40, WL115);
sram_cell_6t_3 inst_cell_115_39 ( BL39, BLN39, WL115);
sram_cell_6t_3 inst_cell_115_38 ( BL38, BLN38, WL115);
sram_cell_6t_3 inst_cell_115_37 ( BL37, BLN37, WL115);
sram_cell_6t_3 inst_cell_115_36 ( BL36, BLN36, WL115);
sram_cell_6t_3 inst_cell_115_35 ( BL35, BLN35, WL115);
sram_cell_6t_3 inst_cell_115_34 ( BL34, BLN34, WL115);
sram_cell_6t_3 inst_cell_115_33 ( BL33, BLN33, WL115);
sram_cell_6t_3 inst_cell_115_32 ( BL32, BLN32, WL115);
sram_cell_6t_3 inst_cell_115_31 ( BL31, BLN31, WL115);
sram_cell_6t_3 inst_cell_115_30 ( BL30, BLN30, WL115);
sram_cell_6t_3 inst_cell_115_29 ( BL29, BLN29, WL115);
sram_cell_6t_3 inst_cell_115_28 ( BL28, BLN28, WL115);
sram_cell_6t_3 inst_cell_115_27 ( BL27, BLN27, WL115);
sram_cell_6t_3 inst_cell_115_26 ( BL26, BLN26, WL115);
sram_cell_6t_3 inst_cell_115_25 ( BL25, BLN25, WL115);
sram_cell_6t_3 inst_cell_115_24 ( BL24, BLN24, WL115);
sram_cell_6t_3 inst_cell_115_23 ( BL23, BLN23, WL115);
sram_cell_6t_3 inst_cell_115_22 ( BL22, BLN22, WL115);
sram_cell_6t_3 inst_cell_115_21 ( BL21, BLN21, WL115);
sram_cell_6t_3 inst_cell_115_20 ( BL20, BLN20, WL115);
sram_cell_6t_3 inst_cell_115_19 ( BL19, BLN19, WL115);
sram_cell_6t_3 inst_cell_115_18 ( BL18, BLN18, WL115);
sram_cell_6t_3 inst_cell_115_17 ( BL17, BLN17, WL115);
sram_cell_6t_3 inst_cell_115_16 ( BL16, BLN16, WL115);
sram_cell_6t_3 inst_cell_115_15 ( BL15, BLN15, WL115);
sram_cell_6t_3 inst_cell_115_14 ( BL14, BLN14, WL115);
sram_cell_6t_3 inst_cell_115_13 ( BL13, BLN13, WL115);
sram_cell_6t_3 inst_cell_115_12 ( BL12, BLN12, WL115);
sram_cell_6t_3 inst_cell_115_11 ( BL11, BLN11, WL115);
sram_cell_6t_3 inst_cell_115_10 ( BL10, BLN10, WL115);
sram_cell_6t_3 inst_cell_115_9 ( BL9, BLN9, WL115);
sram_cell_6t_3 inst_cell_115_8 ( BL8, BLN8, WL115);
sram_cell_6t_3 inst_cell_115_7 ( BL7, BLN7, WL115);
sram_cell_6t_3 inst_cell_115_6 ( BL6, BLN6, WL115);
sram_cell_6t_3 inst_cell_115_5 ( BL5, BLN5, WL115);
sram_cell_6t_3 inst_cell_115_4 ( BL4, BLN4, WL115);
sram_cell_6t_3 inst_cell_115_3 ( BL3, BLN3, WL115);
sram_cell_6t_3 inst_cell_115_2 ( BL2, BLN2, WL115);
sram_cell_6t_3 inst_cell_115_1 ( BL1, BLN1, WL115);
sram_cell_6t_3 inst_cell_115_0 ( BL0, BLN0, WL115);
sram_cell_6t_3 inst_cell_114_127 ( BL127, BLN127, WL114);
sram_cell_6t_3 inst_cell_114_126 ( BL126, BLN126, WL114);
sram_cell_6t_3 inst_cell_114_125 ( BL125, BLN125, WL114);
sram_cell_6t_3 inst_cell_114_124 ( BL124, BLN124, WL114);
sram_cell_6t_3 inst_cell_114_123 ( BL123, BLN123, WL114);
sram_cell_6t_3 inst_cell_114_122 ( BL122, BLN122, WL114);
sram_cell_6t_3 inst_cell_114_121 ( BL121, BLN121, WL114);
sram_cell_6t_3 inst_cell_114_120 ( BL120, BLN120, WL114);
sram_cell_6t_3 inst_cell_114_119 ( BL119, BLN119, WL114);
sram_cell_6t_3 inst_cell_114_118 ( BL118, BLN118, WL114);
sram_cell_6t_3 inst_cell_114_117 ( BL117, BLN117, WL114);
sram_cell_6t_3 inst_cell_114_116 ( BL116, BLN116, WL114);
sram_cell_6t_3 inst_cell_114_115 ( BL115, BLN115, WL114);
sram_cell_6t_3 inst_cell_114_114 ( BL114, BLN114, WL114);
sram_cell_6t_3 inst_cell_114_113 ( BL113, BLN113, WL114);
sram_cell_6t_3 inst_cell_114_112 ( BL112, BLN112, WL114);
sram_cell_6t_3 inst_cell_114_111 ( BL111, BLN111, WL114);
sram_cell_6t_3 inst_cell_114_110 ( BL110, BLN110, WL114);
sram_cell_6t_3 inst_cell_114_109 ( BL109, BLN109, WL114);
sram_cell_6t_3 inst_cell_114_108 ( BL108, BLN108, WL114);
sram_cell_6t_3 inst_cell_114_107 ( BL107, BLN107, WL114);
sram_cell_6t_3 inst_cell_114_106 ( BL106, BLN106, WL114);
sram_cell_6t_3 inst_cell_114_105 ( BL105, BLN105, WL114);
sram_cell_6t_3 inst_cell_114_104 ( BL104, BLN104, WL114);
sram_cell_6t_3 inst_cell_114_103 ( BL103, BLN103, WL114);
sram_cell_6t_3 inst_cell_114_102 ( BL102, BLN102, WL114);
sram_cell_6t_3 inst_cell_114_101 ( BL101, BLN101, WL114);
sram_cell_6t_3 inst_cell_114_100 ( BL100, BLN100, WL114);
sram_cell_6t_3 inst_cell_114_99 ( BL99, BLN99, WL114);
sram_cell_6t_3 inst_cell_114_98 ( BL98, BLN98, WL114);
sram_cell_6t_3 inst_cell_114_97 ( BL97, BLN97, WL114);
sram_cell_6t_3 inst_cell_114_96 ( BL96, BLN96, WL114);
sram_cell_6t_3 inst_cell_114_95 ( BL95, BLN95, WL114);
sram_cell_6t_3 inst_cell_114_94 ( BL94, BLN94, WL114);
sram_cell_6t_3 inst_cell_114_93 ( BL93, BLN93, WL114);
sram_cell_6t_3 inst_cell_114_92 ( BL92, BLN92, WL114);
sram_cell_6t_3 inst_cell_114_91 ( BL91, BLN91, WL114);
sram_cell_6t_3 inst_cell_114_90 ( BL90, BLN90, WL114);
sram_cell_6t_3 inst_cell_114_89 ( BL89, BLN89, WL114);
sram_cell_6t_3 inst_cell_114_88 ( BL88, BLN88, WL114);
sram_cell_6t_3 inst_cell_114_87 ( BL87, BLN87, WL114);
sram_cell_6t_3 inst_cell_114_86 ( BL86, BLN86, WL114);
sram_cell_6t_3 inst_cell_114_85 ( BL85, BLN85, WL114);
sram_cell_6t_3 inst_cell_114_84 ( BL84, BLN84, WL114);
sram_cell_6t_3 inst_cell_114_83 ( BL83, BLN83, WL114);
sram_cell_6t_3 inst_cell_114_82 ( BL82, BLN82, WL114);
sram_cell_6t_3 inst_cell_114_81 ( BL81, BLN81, WL114);
sram_cell_6t_3 inst_cell_114_80 ( BL80, BLN80, WL114);
sram_cell_6t_3 inst_cell_114_79 ( BL79, BLN79, WL114);
sram_cell_6t_3 inst_cell_114_78 ( BL78, BLN78, WL114);
sram_cell_6t_3 inst_cell_114_77 ( BL77, BLN77, WL114);
sram_cell_6t_3 inst_cell_114_76 ( BL76, BLN76, WL114);
sram_cell_6t_3 inst_cell_114_75 ( BL75, BLN75, WL114);
sram_cell_6t_3 inst_cell_114_74 ( BL74, BLN74, WL114);
sram_cell_6t_3 inst_cell_114_73 ( BL73, BLN73, WL114);
sram_cell_6t_3 inst_cell_114_72 ( BL72, BLN72, WL114);
sram_cell_6t_3 inst_cell_114_71 ( BL71, BLN71, WL114);
sram_cell_6t_3 inst_cell_114_70 ( BL70, BLN70, WL114);
sram_cell_6t_3 inst_cell_114_69 ( BL69, BLN69, WL114);
sram_cell_6t_3 inst_cell_114_68 ( BL68, BLN68, WL114);
sram_cell_6t_3 inst_cell_114_67 ( BL67, BLN67, WL114);
sram_cell_6t_3 inst_cell_114_66 ( BL66, BLN66, WL114);
sram_cell_6t_3 inst_cell_114_65 ( BL65, BLN65, WL114);
sram_cell_6t_3 inst_cell_114_64 ( BL64, BLN64, WL114);
sram_cell_6t_3 inst_cell_114_63 ( BL63, BLN63, WL114);
sram_cell_6t_3 inst_cell_114_62 ( BL62, BLN62, WL114);
sram_cell_6t_3 inst_cell_114_61 ( BL61, BLN61, WL114);
sram_cell_6t_3 inst_cell_114_60 ( BL60, BLN60, WL114);
sram_cell_6t_3 inst_cell_114_59 ( BL59, BLN59, WL114);
sram_cell_6t_3 inst_cell_114_58 ( BL58, BLN58, WL114);
sram_cell_6t_3 inst_cell_114_57 ( BL57, BLN57, WL114);
sram_cell_6t_3 inst_cell_114_56 ( BL56, BLN56, WL114);
sram_cell_6t_3 inst_cell_114_55 ( BL55, BLN55, WL114);
sram_cell_6t_3 inst_cell_114_54 ( BL54, BLN54, WL114);
sram_cell_6t_3 inst_cell_114_53 ( BL53, BLN53, WL114);
sram_cell_6t_3 inst_cell_114_52 ( BL52, BLN52, WL114);
sram_cell_6t_3 inst_cell_114_51 ( BL51, BLN51, WL114);
sram_cell_6t_3 inst_cell_114_50 ( BL50, BLN50, WL114);
sram_cell_6t_3 inst_cell_114_49 ( BL49, BLN49, WL114);
sram_cell_6t_3 inst_cell_114_48 ( BL48, BLN48, WL114);
sram_cell_6t_3 inst_cell_114_47 ( BL47, BLN47, WL114);
sram_cell_6t_3 inst_cell_114_46 ( BL46, BLN46, WL114);
sram_cell_6t_3 inst_cell_114_45 ( BL45, BLN45, WL114);
sram_cell_6t_3 inst_cell_114_44 ( BL44, BLN44, WL114);
sram_cell_6t_3 inst_cell_114_43 ( BL43, BLN43, WL114);
sram_cell_6t_3 inst_cell_114_42 ( BL42, BLN42, WL114);
sram_cell_6t_3 inst_cell_114_41 ( BL41, BLN41, WL114);
sram_cell_6t_3 inst_cell_114_40 ( BL40, BLN40, WL114);
sram_cell_6t_3 inst_cell_114_39 ( BL39, BLN39, WL114);
sram_cell_6t_3 inst_cell_114_38 ( BL38, BLN38, WL114);
sram_cell_6t_3 inst_cell_114_37 ( BL37, BLN37, WL114);
sram_cell_6t_3 inst_cell_114_36 ( BL36, BLN36, WL114);
sram_cell_6t_3 inst_cell_114_35 ( BL35, BLN35, WL114);
sram_cell_6t_3 inst_cell_114_34 ( BL34, BLN34, WL114);
sram_cell_6t_3 inst_cell_114_33 ( BL33, BLN33, WL114);
sram_cell_6t_3 inst_cell_114_32 ( BL32, BLN32, WL114);
sram_cell_6t_3 inst_cell_114_31 ( BL31, BLN31, WL114);
sram_cell_6t_3 inst_cell_114_30 ( BL30, BLN30, WL114);
sram_cell_6t_3 inst_cell_114_29 ( BL29, BLN29, WL114);
sram_cell_6t_3 inst_cell_114_28 ( BL28, BLN28, WL114);
sram_cell_6t_3 inst_cell_114_27 ( BL27, BLN27, WL114);
sram_cell_6t_3 inst_cell_114_26 ( BL26, BLN26, WL114);
sram_cell_6t_3 inst_cell_114_25 ( BL25, BLN25, WL114);
sram_cell_6t_3 inst_cell_114_24 ( BL24, BLN24, WL114);
sram_cell_6t_3 inst_cell_114_23 ( BL23, BLN23, WL114);
sram_cell_6t_3 inst_cell_114_22 ( BL22, BLN22, WL114);
sram_cell_6t_3 inst_cell_114_21 ( BL21, BLN21, WL114);
sram_cell_6t_3 inst_cell_114_20 ( BL20, BLN20, WL114);
sram_cell_6t_3 inst_cell_114_19 ( BL19, BLN19, WL114);
sram_cell_6t_3 inst_cell_114_18 ( BL18, BLN18, WL114);
sram_cell_6t_3 inst_cell_114_17 ( BL17, BLN17, WL114);
sram_cell_6t_3 inst_cell_114_16 ( BL16, BLN16, WL114);
sram_cell_6t_3 inst_cell_114_15 ( BL15, BLN15, WL114);
sram_cell_6t_3 inst_cell_114_14 ( BL14, BLN14, WL114);
sram_cell_6t_3 inst_cell_114_13 ( BL13, BLN13, WL114);
sram_cell_6t_3 inst_cell_114_12 ( BL12, BLN12, WL114);
sram_cell_6t_3 inst_cell_114_11 ( BL11, BLN11, WL114);
sram_cell_6t_3 inst_cell_114_10 ( BL10, BLN10, WL114);
sram_cell_6t_3 inst_cell_114_9 ( BL9, BLN9, WL114);
sram_cell_6t_3 inst_cell_114_8 ( BL8, BLN8, WL114);
sram_cell_6t_3 inst_cell_114_7 ( BL7, BLN7, WL114);
sram_cell_6t_3 inst_cell_114_6 ( BL6, BLN6, WL114);
sram_cell_6t_3 inst_cell_114_5 ( BL5, BLN5, WL114);
sram_cell_6t_3 inst_cell_114_4 ( BL4, BLN4, WL114);
sram_cell_6t_3 inst_cell_114_3 ( BL3, BLN3, WL114);
sram_cell_6t_3 inst_cell_114_2 ( BL2, BLN2, WL114);
sram_cell_6t_3 inst_cell_114_1 ( BL1, BLN1, WL114);
sram_cell_6t_3 inst_cell_114_0 ( BL0, BLN0, WL114);
sram_cell_6t_3 inst_cell_113_127 ( BL127, BLN127, WL113);
sram_cell_6t_3 inst_cell_113_126 ( BL126, BLN126, WL113);
sram_cell_6t_3 inst_cell_113_125 ( BL125, BLN125, WL113);
sram_cell_6t_3 inst_cell_113_124 ( BL124, BLN124, WL113);
sram_cell_6t_3 inst_cell_113_123 ( BL123, BLN123, WL113);
sram_cell_6t_3 inst_cell_113_122 ( BL122, BLN122, WL113);
sram_cell_6t_3 inst_cell_113_121 ( BL121, BLN121, WL113);
sram_cell_6t_3 inst_cell_113_120 ( BL120, BLN120, WL113);
sram_cell_6t_3 inst_cell_113_119 ( BL119, BLN119, WL113);
sram_cell_6t_3 inst_cell_113_118 ( BL118, BLN118, WL113);
sram_cell_6t_3 inst_cell_113_117 ( BL117, BLN117, WL113);
sram_cell_6t_3 inst_cell_113_116 ( BL116, BLN116, WL113);
sram_cell_6t_3 inst_cell_113_115 ( BL115, BLN115, WL113);
sram_cell_6t_3 inst_cell_113_114 ( BL114, BLN114, WL113);
sram_cell_6t_3 inst_cell_113_113 ( BL113, BLN113, WL113);
sram_cell_6t_3 inst_cell_113_112 ( BL112, BLN112, WL113);
sram_cell_6t_3 inst_cell_113_111 ( BL111, BLN111, WL113);
sram_cell_6t_3 inst_cell_113_110 ( BL110, BLN110, WL113);
sram_cell_6t_3 inst_cell_113_109 ( BL109, BLN109, WL113);
sram_cell_6t_3 inst_cell_113_108 ( BL108, BLN108, WL113);
sram_cell_6t_3 inst_cell_113_107 ( BL107, BLN107, WL113);
sram_cell_6t_3 inst_cell_113_106 ( BL106, BLN106, WL113);
sram_cell_6t_3 inst_cell_113_105 ( BL105, BLN105, WL113);
sram_cell_6t_3 inst_cell_113_104 ( BL104, BLN104, WL113);
sram_cell_6t_3 inst_cell_113_103 ( BL103, BLN103, WL113);
sram_cell_6t_3 inst_cell_113_102 ( BL102, BLN102, WL113);
sram_cell_6t_3 inst_cell_113_101 ( BL101, BLN101, WL113);
sram_cell_6t_3 inst_cell_113_100 ( BL100, BLN100, WL113);
sram_cell_6t_3 inst_cell_113_99 ( BL99, BLN99, WL113);
sram_cell_6t_3 inst_cell_113_98 ( BL98, BLN98, WL113);
sram_cell_6t_3 inst_cell_113_97 ( BL97, BLN97, WL113);
sram_cell_6t_3 inst_cell_113_96 ( BL96, BLN96, WL113);
sram_cell_6t_3 inst_cell_113_95 ( BL95, BLN95, WL113);
sram_cell_6t_3 inst_cell_113_94 ( BL94, BLN94, WL113);
sram_cell_6t_3 inst_cell_113_93 ( BL93, BLN93, WL113);
sram_cell_6t_3 inst_cell_113_92 ( BL92, BLN92, WL113);
sram_cell_6t_3 inst_cell_113_91 ( BL91, BLN91, WL113);
sram_cell_6t_3 inst_cell_113_90 ( BL90, BLN90, WL113);
sram_cell_6t_3 inst_cell_113_89 ( BL89, BLN89, WL113);
sram_cell_6t_3 inst_cell_113_88 ( BL88, BLN88, WL113);
sram_cell_6t_3 inst_cell_113_87 ( BL87, BLN87, WL113);
sram_cell_6t_3 inst_cell_113_86 ( BL86, BLN86, WL113);
sram_cell_6t_3 inst_cell_113_85 ( BL85, BLN85, WL113);
sram_cell_6t_3 inst_cell_113_84 ( BL84, BLN84, WL113);
sram_cell_6t_3 inst_cell_113_83 ( BL83, BLN83, WL113);
sram_cell_6t_3 inst_cell_113_82 ( BL82, BLN82, WL113);
sram_cell_6t_3 inst_cell_113_81 ( BL81, BLN81, WL113);
sram_cell_6t_3 inst_cell_113_80 ( BL80, BLN80, WL113);
sram_cell_6t_3 inst_cell_113_79 ( BL79, BLN79, WL113);
sram_cell_6t_3 inst_cell_113_78 ( BL78, BLN78, WL113);
sram_cell_6t_3 inst_cell_113_77 ( BL77, BLN77, WL113);
sram_cell_6t_3 inst_cell_113_76 ( BL76, BLN76, WL113);
sram_cell_6t_3 inst_cell_113_75 ( BL75, BLN75, WL113);
sram_cell_6t_3 inst_cell_113_74 ( BL74, BLN74, WL113);
sram_cell_6t_3 inst_cell_113_73 ( BL73, BLN73, WL113);
sram_cell_6t_3 inst_cell_113_72 ( BL72, BLN72, WL113);
sram_cell_6t_3 inst_cell_113_71 ( BL71, BLN71, WL113);
sram_cell_6t_3 inst_cell_113_70 ( BL70, BLN70, WL113);
sram_cell_6t_3 inst_cell_113_69 ( BL69, BLN69, WL113);
sram_cell_6t_3 inst_cell_113_68 ( BL68, BLN68, WL113);
sram_cell_6t_3 inst_cell_113_67 ( BL67, BLN67, WL113);
sram_cell_6t_3 inst_cell_113_66 ( BL66, BLN66, WL113);
sram_cell_6t_3 inst_cell_113_65 ( BL65, BLN65, WL113);
sram_cell_6t_3 inst_cell_113_64 ( BL64, BLN64, WL113);
sram_cell_6t_3 inst_cell_113_63 ( BL63, BLN63, WL113);
sram_cell_6t_3 inst_cell_113_62 ( BL62, BLN62, WL113);
sram_cell_6t_3 inst_cell_113_61 ( BL61, BLN61, WL113);
sram_cell_6t_3 inst_cell_113_60 ( BL60, BLN60, WL113);
sram_cell_6t_3 inst_cell_113_59 ( BL59, BLN59, WL113);
sram_cell_6t_3 inst_cell_113_58 ( BL58, BLN58, WL113);
sram_cell_6t_3 inst_cell_113_57 ( BL57, BLN57, WL113);
sram_cell_6t_3 inst_cell_113_56 ( BL56, BLN56, WL113);
sram_cell_6t_3 inst_cell_113_55 ( BL55, BLN55, WL113);
sram_cell_6t_3 inst_cell_113_54 ( BL54, BLN54, WL113);
sram_cell_6t_3 inst_cell_113_53 ( BL53, BLN53, WL113);
sram_cell_6t_3 inst_cell_113_52 ( BL52, BLN52, WL113);
sram_cell_6t_3 inst_cell_113_51 ( BL51, BLN51, WL113);
sram_cell_6t_3 inst_cell_113_50 ( BL50, BLN50, WL113);
sram_cell_6t_3 inst_cell_113_49 ( BL49, BLN49, WL113);
sram_cell_6t_3 inst_cell_113_48 ( BL48, BLN48, WL113);
sram_cell_6t_3 inst_cell_113_47 ( BL47, BLN47, WL113);
sram_cell_6t_3 inst_cell_113_46 ( BL46, BLN46, WL113);
sram_cell_6t_3 inst_cell_113_45 ( BL45, BLN45, WL113);
sram_cell_6t_3 inst_cell_113_44 ( BL44, BLN44, WL113);
sram_cell_6t_3 inst_cell_113_43 ( BL43, BLN43, WL113);
sram_cell_6t_3 inst_cell_113_42 ( BL42, BLN42, WL113);
sram_cell_6t_3 inst_cell_113_41 ( BL41, BLN41, WL113);
sram_cell_6t_3 inst_cell_113_40 ( BL40, BLN40, WL113);
sram_cell_6t_3 inst_cell_113_39 ( BL39, BLN39, WL113);
sram_cell_6t_3 inst_cell_113_38 ( BL38, BLN38, WL113);
sram_cell_6t_3 inst_cell_113_37 ( BL37, BLN37, WL113);
sram_cell_6t_3 inst_cell_113_36 ( BL36, BLN36, WL113);
sram_cell_6t_3 inst_cell_113_35 ( BL35, BLN35, WL113);
sram_cell_6t_3 inst_cell_113_34 ( BL34, BLN34, WL113);
sram_cell_6t_3 inst_cell_113_33 ( BL33, BLN33, WL113);
sram_cell_6t_3 inst_cell_113_32 ( BL32, BLN32, WL113);
sram_cell_6t_3 inst_cell_113_31 ( BL31, BLN31, WL113);
sram_cell_6t_3 inst_cell_113_30 ( BL30, BLN30, WL113);
sram_cell_6t_3 inst_cell_113_29 ( BL29, BLN29, WL113);
sram_cell_6t_3 inst_cell_113_28 ( BL28, BLN28, WL113);
sram_cell_6t_3 inst_cell_113_27 ( BL27, BLN27, WL113);
sram_cell_6t_3 inst_cell_113_26 ( BL26, BLN26, WL113);
sram_cell_6t_3 inst_cell_113_25 ( BL25, BLN25, WL113);
sram_cell_6t_3 inst_cell_113_24 ( BL24, BLN24, WL113);
sram_cell_6t_3 inst_cell_113_23 ( BL23, BLN23, WL113);
sram_cell_6t_3 inst_cell_113_22 ( BL22, BLN22, WL113);
sram_cell_6t_3 inst_cell_113_21 ( BL21, BLN21, WL113);
sram_cell_6t_3 inst_cell_113_20 ( BL20, BLN20, WL113);
sram_cell_6t_3 inst_cell_113_19 ( BL19, BLN19, WL113);
sram_cell_6t_3 inst_cell_113_18 ( BL18, BLN18, WL113);
sram_cell_6t_3 inst_cell_113_17 ( BL17, BLN17, WL113);
sram_cell_6t_3 inst_cell_113_16 ( BL16, BLN16, WL113);
sram_cell_6t_3 inst_cell_113_15 ( BL15, BLN15, WL113);
sram_cell_6t_3 inst_cell_113_14 ( BL14, BLN14, WL113);
sram_cell_6t_3 inst_cell_113_13 ( BL13, BLN13, WL113);
sram_cell_6t_3 inst_cell_113_12 ( BL12, BLN12, WL113);
sram_cell_6t_3 inst_cell_113_11 ( BL11, BLN11, WL113);
sram_cell_6t_3 inst_cell_113_10 ( BL10, BLN10, WL113);
sram_cell_6t_3 inst_cell_113_9 ( BL9, BLN9, WL113);
sram_cell_6t_3 inst_cell_113_8 ( BL8, BLN8, WL113);
sram_cell_6t_3 inst_cell_113_7 ( BL7, BLN7, WL113);
sram_cell_6t_3 inst_cell_113_6 ( BL6, BLN6, WL113);
sram_cell_6t_3 inst_cell_113_5 ( BL5, BLN5, WL113);
sram_cell_6t_3 inst_cell_113_4 ( BL4, BLN4, WL113);
sram_cell_6t_3 inst_cell_113_3 ( BL3, BLN3, WL113);
sram_cell_6t_3 inst_cell_113_2 ( BL2, BLN2, WL113);
sram_cell_6t_3 inst_cell_113_1 ( BL1, BLN1, WL113);
sram_cell_6t_3 inst_cell_113_0 ( BL0, BLN0, WL113);
sram_cell_6t_3 inst_cell_112_127 ( BL127, BLN127, WL112);
sram_cell_6t_3 inst_cell_112_126 ( BL126, BLN126, WL112);
sram_cell_6t_3 inst_cell_112_125 ( BL125, BLN125, WL112);
sram_cell_6t_3 inst_cell_112_124 ( BL124, BLN124, WL112);
sram_cell_6t_3 inst_cell_112_123 ( BL123, BLN123, WL112);
sram_cell_6t_3 inst_cell_112_122 ( BL122, BLN122, WL112);
sram_cell_6t_3 inst_cell_112_121 ( BL121, BLN121, WL112);
sram_cell_6t_3 inst_cell_112_120 ( BL120, BLN120, WL112);
sram_cell_6t_3 inst_cell_112_119 ( BL119, BLN119, WL112);
sram_cell_6t_3 inst_cell_112_118 ( BL118, BLN118, WL112);
sram_cell_6t_3 inst_cell_112_117 ( BL117, BLN117, WL112);
sram_cell_6t_3 inst_cell_112_116 ( BL116, BLN116, WL112);
sram_cell_6t_3 inst_cell_112_115 ( BL115, BLN115, WL112);
sram_cell_6t_3 inst_cell_112_114 ( BL114, BLN114, WL112);
sram_cell_6t_3 inst_cell_112_113 ( BL113, BLN113, WL112);
sram_cell_6t_3 inst_cell_112_112 ( BL112, BLN112, WL112);
sram_cell_6t_3 inst_cell_112_111 ( BL111, BLN111, WL112);
sram_cell_6t_3 inst_cell_112_110 ( BL110, BLN110, WL112);
sram_cell_6t_3 inst_cell_112_109 ( BL109, BLN109, WL112);
sram_cell_6t_3 inst_cell_112_108 ( BL108, BLN108, WL112);
sram_cell_6t_3 inst_cell_112_107 ( BL107, BLN107, WL112);
sram_cell_6t_3 inst_cell_112_106 ( BL106, BLN106, WL112);
sram_cell_6t_3 inst_cell_112_105 ( BL105, BLN105, WL112);
sram_cell_6t_3 inst_cell_112_104 ( BL104, BLN104, WL112);
sram_cell_6t_3 inst_cell_112_103 ( BL103, BLN103, WL112);
sram_cell_6t_3 inst_cell_112_102 ( BL102, BLN102, WL112);
sram_cell_6t_3 inst_cell_112_101 ( BL101, BLN101, WL112);
sram_cell_6t_3 inst_cell_112_100 ( BL100, BLN100, WL112);
sram_cell_6t_3 inst_cell_112_99 ( BL99, BLN99, WL112);
sram_cell_6t_3 inst_cell_112_98 ( BL98, BLN98, WL112);
sram_cell_6t_3 inst_cell_112_97 ( BL97, BLN97, WL112);
sram_cell_6t_3 inst_cell_112_96 ( BL96, BLN96, WL112);
sram_cell_6t_3 inst_cell_112_95 ( BL95, BLN95, WL112);
sram_cell_6t_3 inst_cell_112_94 ( BL94, BLN94, WL112);
sram_cell_6t_3 inst_cell_112_93 ( BL93, BLN93, WL112);
sram_cell_6t_3 inst_cell_112_92 ( BL92, BLN92, WL112);
sram_cell_6t_3 inst_cell_112_91 ( BL91, BLN91, WL112);
sram_cell_6t_3 inst_cell_112_90 ( BL90, BLN90, WL112);
sram_cell_6t_3 inst_cell_112_89 ( BL89, BLN89, WL112);
sram_cell_6t_3 inst_cell_112_88 ( BL88, BLN88, WL112);
sram_cell_6t_3 inst_cell_112_87 ( BL87, BLN87, WL112);
sram_cell_6t_3 inst_cell_112_86 ( BL86, BLN86, WL112);
sram_cell_6t_3 inst_cell_112_85 ( BL85, BLN85, WL112);
sram_cell_6t_3 inst_cell_112_84 ( BL84, BLN84, WL112);
sram_cell_6t_3 inst_cell_112_83 ( BL83, BLN83, WL112);
sram_cell_6t_3 inst_cell_112_82 ( BL82, BLN82, WL112);
sram_cell_6t_3 inst_cell_112_81 ( BL81, BLN81, WL112);
sram_cell_6t_3 inst_cell_112_80 ( BL80, BLN80, WL112);
sram_cell_6t_3 inst_cell_112_79 ( BL79, BLN79, WL112);
sram_cell_6t_3 inst_cell_112_78 ( BL78, BLN78, WL112);
sram_cell_6t_3 inst_cell_112_77 ( BL77, BLN77, WL112);
sram_cell_6t_3 inst_cell_112_76 ( BL76, BLN76, WL112);
sram_cell_6t_3 inst_cell_112_75 ( BL75, BLN75, WL112);
sram_cell_6t_3 inst_cell_112_74 ( BL74, BLN74, WL112);
sram_cell_6t_3 inst_cell_112_73 ( BL73, BLN73, WL112);
sram_cell_6t_3 inst_cell_112_72 ( BL72, BLN72, WL112);
sram_cell_6t_3 inst_cell_112_71 ( BL71, BLN71, WL112);
sram_cell_6t_3 inst_cell_112_70 ( BL70, BLN70, WL112);
sram_cell_6t_3 inst_cell_112_69 ( BL69, BLN69, WL112);
sram_cell_6t_3 inst_cell_112_68 ( BL68, BLN68, WL112);
sram_cell_6t_3 inst_cell_112_67 ( BL67, BLN67, WL112);
sram_cell_6t_3 inst_cell_112_66 ( BL66, BLN66, WL112);
sram_cell_6t_3 inst_cell_112_65 ( BL65, BLN65, WL112);
sram_cell_6t_3 inst_cell_112_64 ( BL64, BLN64, WL112);
sram_cell_6t_3 inst_cell_112_63 ( BL63, BLN63, WL112);
sram_cell_6t_3 inst_cell_112_62 ( BL62, BLN62, WL112);
sram_cell_6t_3 inst_cell_112_61 ( BL61, BLN61, WL112);
sram_cell_6t_3 inst_cell_112_60 ( BL60, BLN60, WL112);
sram_cell_6t_3 inst_cell_112_59 ( BL59, BLN59, WL112);
sram_cell_6t_3 inst_cell_112_58 ( BL58, BLN58, WL112);
sram_cell_6t_3 inst_cell_112_57 ( BL57, BLN57, WL112);
sram_cell_6t_3 inst_cell_112_56 ( BL56, BLN56, WL112);
sram_cell_6t_3 inst_cell_112_55 ( BL55, BLN55, WL112);
sram_cell_6t_3 inst_cell_112_54 ( BL54, BLN54, WL112);
sram_cell_6t_3 inst_cell_112_53 ( BL53, BLN53, WL112);
sram_cell_6t_3 inst_cell_112_52 ( BL52, BLN52, WL112);
sram_cell_6t_3 inst_cell_112_51 ( BL51, BLN51, WL112);
sram_cell_6t_3 inst_cell_112_50 ( BL50, BLN50, WL112);
sram_cell_6t_3 inst_cell_112_49 ( BL49, BLN49, WL112);
sram_cell_6t_3 inst_cell_112_48 ( BL48, BLN48, WL112);
sram_cell_6t_3 inst_cell_112_47 ( BL47, BLN47, WL112);
sram_cell_6t_3 inst_cell_112_46 ( BL46, BLN46, WL112);
sram_cell_6t_3 inst_cell_112_45 ( BL45, BLN45, WL112);
sram_cell_6t_3 inst_cell_112_44 ( BL44, BLN44, WL112);
sram_cell_6t_3 inst_cell_112_43 ( BL43, BLN43, WL112);
sram_cell_6t_3 inst_cell_112_42 ( BL42, BLN42, WL112);
sram_cell_6t_3 inst_cell_112_41 ( BL41, BLN41, WL112);
sram_cell_6t_3 inst_cell_112_40 ( BL40, BLN40, WL112);
sram_cell_6t_3 inst_cell_112_39 ( BL39, BLN39, WL112);
sram_cell_6t_3 inst_cell_112_38 ( BL38, BLN38, WL112);
sram_cell_6t_3 inst_cell_112_37 ( BL37, BLN37, WL112);
sram_cell_6t_3 inst_cell_112_36 ( BL36, BLN36, WL112);
sram_cell_6t_3 inst_cell_112_35 ( BL35, BLN35, WL112);
sram_cell_6t_3 inst_cell_112_34 ( BL34, BLN34, WL112);
sram_cell_6t_3 inst_cell_112_33 ( BL33, BLN33, WL112);
sram_cell_6t_3 inst_cell_112_32 ( BL32, BLN32, WL112);
sram_cell_6t_3 inst_cell_112_31 ( BL31, BLN31, WL112);
sram_cell_6t_3 inst_cell_112_30 ( BL30, BLN30, WL112);
sram_cell_6t_3 inst_cell_112_29 ( BL29, BLN29, WL112);
sram_cell_6t_3 inst_cell_112_28 ( BL28, BLN28, WL112);
sram_cell_6t_3 inst_cell_112_27 ( BL27, BLN27, WL112);
sram_cell_6t_3 inst_cell_112_26 ( BL26, BLN26, WL112);
sram_cell_6t_3 inst_cell_112_25 ( BL25, BLN25, WL112);
sram_cell_6t_3 inst_cell_112_24 ( BL24, BLN24, WL112);
sram_cell_6t_3 inst_cell_112_23 ( BL23, BLN23, WL112);
sram_cell_6t_3 inst_cell_112_22 ( BL22, BLN22, WL112);
sram_cell_6t_3 inst_cell_112_21 ( BL21, BLN21, WL112);
sram_cell_6t_3 inst_cell_112_20 ( BL20, BLN20, WL112);
sram_cell_6t_3 inst_cell_112_19 ( BL19, BLN19, WL112);
sram_cell_6t_3 inst_cell_112_18 ( BL18, BLN18, WL112);
sram_cell_6t_3 inst_cell_112_17 ( BL17, BLN17, WL112);
sram_cell_6t_3 inst_cell_112_16 ( BL16, BLN16, WL112);
sram_cell_6t_3 inst_cell_112_15 ( BL15, BLN15, WL112);
sram_cell_6t_3 inst_cell_112_14 ( BL14, BLN14, WL112);
sram_cell_6t_3 inst_cell_112_13 ( BL13, BLN13, WL112);
sram_cell_6t_3 inst_cell_112_12 ( BL12, BLN12, WL112);
sram_cell_6t_3 inst_cell_112_11 ( BL11, BLN11, WL112);
sram_cell_6t_3 inst_cell_112_10 ( BL10, BLN10, WL112);
sram_cell_6t_3 inst_cell_112_9 ( BL9, BLN9, WL112);
sram_cell_6t_3 inst_cell_112_8 ( BL8, BLN8, WL112);
sram_cell_6t_3 inst_cell_112_7 ( BL7, BLN7, WL112);
sram_cell_6t_3 inst_cell_112_6 ( BL6, BLN6, WL112);
sram_cell_6t_3 inst_cell_112_5 ( BL5, BLN5, WL112);
sram_cell_6t_3 inst_cell_112_4 ( BL4, BLN4, WL112);
sram_cell_6t_3 inst_cell_112_3 ( BL3, BLN3, WL112);
sram_cell_6t_3 inst_cell_112_2 ( BL2, BLN2, WL112);
sram_cell_6t_3 inst_cell_112_1 ( BL1, BLN1, WL112);
sram_cell_6t_3 inst_cell_112_0 ( BL0, BLN0, WL112);
sram_cell_6t_3 inst_cell_111_127 ( BL127, BLN127, WL111);
sram_cell_6t_3 inst_cell_111_126 ( BL126, BLN126, WL111);
sram_cell_6t_3 inst_cell_111_125 ( BL125, BLN125, WL111);
sram_cell_6t_3 inst_cell_111_124 ( BL124, BLN124, WL111);
sram_cell_6t_3 inst_cell_111_123 ( BL123, BLN123, WL111);
sram_cell_6t_3 inst_cell_111_122 ( BL122, BLN122, WL111);
sram_cell_6t_3 inst_cell_111_121 ( BL121, BLN121, WL111);
sram_cell_6t_3 inst_cell_111_120 ( BL120, BLN120, WL111);
sram_cell_6t_3 inst_cell_111_119 ( BL119, BLN119, WL111);
sram_cell_6t_3 inst_cell_111_118 ( BL118, BLN118, WL111);
sram_cell_6t_3 inst_cell_111_117 ( BL117, BLN117, WL111);
sram_cell_6t_3 inst_cell_111_116 ( BL116, BLN116, WL111);
sram_cell_6t_3 inst_cell_111_115 ( BL115, BLN115, WL111);
sram_cell_6t_3 inst_cell_111_114 ( BL114, BLN114, WL111);
sram_cell_6t_3 inst_cell_111_113 ( BL113, BLN113, WL111);
sram_cell_6t_3 inst_cell_111_112 ( BL112, BLN112, WL111);
sram_cell_6t_3 inst_cell_111_111 ( BL111, BLN111, WL111);
sram_cell_6t_3 inst_cell_111_110 ( BL110, BLN110, WL111);
sram_cell_6t_3 inst_cell_111_109 ( BL109, BLN109, WL111);
sram_cell_6t_3 inst_cell_111_108 ( BL108, BLN108, WL111);
sram_cell_6t_3 inst_cell_111_107 ( BL107, BLN107, WL111);
sram_cell_6t_3 inst_cell_111_106 ( BL106, BLN106, WL111);
sram_cell_6t_3 inst_cell_111_105 ( BL105, BLN105, WL111);
sram_cell_6t_3 inst_cell_111_104 ( BL104, BLN104, WL111);
sram_cell_6t_3 inst_cell_111_103 ( BL103, BLN103, WL111);
sram_cell_6t_3 inst_cell_111_102 ( BL102, BLN102, WL111);
sram_cell_6t_3 inst_cell_111_101 ( BL101, BLN101, WL111);
sram_cell_6t_3 inst_cell_111_100 ( BL100, BLN100, WL111);
sram_cell_6t_3 inst_cell_111_99 ( BL99, BLN99, WL111);
sram_cell_6t_3 inst_cell_111_98 ( BL98, BLN98, WL111);
sram_cell_6t_3 inst_cell_111_97 ( BL97, BLN97, WL111);
sram_cell_6t_3 inst_cell_111_96 ( BL96, BLN96, WL111);
sram_cell_6t_3 inst_cell_111_95 ( BL95, BLN95, WL111);
sram_cell_6t_3 inst_cell_111_94 ( BL94, BLN94, WL111);
sram_cell_6t_3 inst_cell_111_93 ( BL93, BLN93, WL111);
sram_cell_6t_3 inst_cell_111_92 ( BL92, BLN92, WL111);
sram_cell_6t_3 inst_cell_111_91 ( BL91, BLN91, WL111);
sram_cell_6t_3 inst_cell_111_90 ( BL90, BLN90, WL111);
sram_cell_6t_3 inst_cell_111_89 ( BL89, BLN89, WL111);
sram_cell_6t_3 inst_cell_111_88 ( BL88, BLN88, WL111);
sram_cell_6t_3 inst_cell_111_87 ( BL87, BLN87, WL111);
sram_cell_6t_3 inst_cell_111_86 ( BL86, BLN86, WL111);
sram_cell_6t_3 inst_cell_111_85 ( BL85, BLN85, WL111);
sram_cell_6t_3 inst_cell_111_84 ( BL84, BLN84, WL111);
sram_cell_6t_3 inst_cell_111_83 ( BL83, BLN83, WL111);
sram_cell_6t_3 inst_cell_111_82 ( BL82, BLN82, WL111);
sram_cell_6t_3 inst_cell_111_81 ( BL81, BLN81, WL111);
sram_cell_6t_3 inst_cell_111_80 ( BL80, BLN80, WL111);
sram_cell_6t_3 inst_cell_111_79 ( BL79, BLN79, WL111);
sram_cell_6t_3 inst_cell_111_78 ( BL78, BLN78, WL111);
sram_cell_6t_3 inst_cell_111_77 ( BL77, BLN77, WL111);
sram_cell_6t_3 inst_cell_111_76 ( BL76, BLN76, WL111);
sram_cell_6t_3 inst_cell_111_75 ( BL75, BLN75, WL111);
sram_cell_6t_3 inst_cell_111_74 ( BL74, BLN74, WL111);
sram_cell_6t_3 inst_cell_111_73 ( BL73, BLN73, WL111);
sram_cell_6t_3 inst_cell_111_72 ( BL72, BLN72, WL111);
sram_cell_6t_3 inst_cell_111_71 ( BL71, BLN71, WL111);
sram_cell_6t_3 inst_cell_111_70 ( BL70, BLN70, WL111);
sram_cell_6t_3 inst_cell_111_69 ( BL69, BLN69, WL111);
sram_cell_6t_3 inst_cell_111_68 ( BL68, BLN68, WL111);
sram_cell_6t_3 inst_cell_111_67 ( BL67, BLN67, WL111);
sram_cell_6t_3 inst_cell_111_66 ( BL66, BLN66, WL111);
sram_cell_6t_3 inst_cell_111_65 ( BL65, BLN65, WL111);
sram_cell_6t_3 inst_cell_111_64 ( BL64, BLN64, WL111);
sram_cell_6t_3 inst_cell_111_63 ( BL63, BLN63, WL111);
sram_cell_6t_3 inst_cell_111_62 ( BL62, BLN62, WL111);
sram_cell_6t_3 inst_cell_111_61 ( BL61, BLN61, WL111);
sram_cell_6t_3 inst_cell_111_60 ( BL60, BLN60, WL111);
sram_cell_6t_3 inst_cell_111_59 ( BL59, BLN59, WL111);
sram_cell_6t_3 inst_cell_111_58 ( BL58, BLN58, WL111);
sram_cell_6t_3 inst_cell_111_57 ( BL57, BLN57, WL111);
sram_cell_6t_3 inst_cell_111_56 ( BL56, BLN56, WL111);
sram_cell_6t_3 inst_cell_111_55 ( BL55, BLN55, WL111);
sram_cell_6t_3 inst_cell_111_54 ( BL54, BLN54, WL111);
sram_cell_6t_3 inst_cell_111_53 ( BL53, BLN53, WL111);
sram_cell_6t_3 inst_cell_111_52 ( BL52, BLN52, WL111);
sram_cell_6t_3 inst_cell_111_51 ( BL51, BLN51, WL111);
sram_cell_6t_3 inst_cell_111_50 ( BL50, BLN50, WL111);
sram_cell_6t_3 inst_cell_111_49 ( BL49, BLN49, WL111);
sram_cell_6t_3 inst_cell_111_48 ( BL48, BLN48, WL111);
sram_cell_6t_3 inst_cell_111_47 ( BL47, BLN47, WL111);
sram_cell_6t_3 inst_cell_111_46 ( BL46, BLN46, WL111);
sram_cell_6t_3 inst_cell_111_45 ( BL45, BLN45, WL111);
sram_cell_6t_3 inst_cell_111_44 ( BL44, BLN44, WL111);
sram_cell_6t_3 inst_cell_111_43 ( BL43, BLN43, WL111);
sram_cell_6t_3 inst_cell_111_42 ( BL42, BLN42, WL111);
sram_cell_6t_3 inst_cell_111_41 ( BL41, BLN41, WL111);
sram_cell_6t_3 inst_cell_111_40 ( BL40, BLN40, WL111);
sram_cell_6t_3 inst_cell_111_39 ( BL39, BLN39, WL111);
sram_cell_6t_3 inst_cell_111_38 ( BL38, BLN38, WL111);
sram_cell_6t_3 inst_cell_111_37 ( BL37, BLN37, WL111);
sram_cell_6t_3 inst_cell_111_36 ( BL36, BLN36, WL111);
sram_cell_6t_3 inst_cell_111_35 ( BL35, BLN35, WL111);
sram_cell_6t_3 inst_cell_111_34 ( BL34, BLN34, WL111);
sram_cell_6t_3 inst_cell_111_33 ( BL33, BLN33, WL111);
sram_cell_6t_3 inst_cell_111_32 ( BL32, BLN32, WL111);
sram_cell_6t_3 inst_cell_111_31 ( BL31, BLN31, WL111);
sram_cell_6t_3 inst_cell_111_30 ( BL30, BLN30, WL111);
sram_cell_6t_3 inst_cell_111_29 ( BL29, BLN29, WL111);
sram_cell_6t_3 inst_cell_111_28 ( BL28, BLN28, WL111);
sram_cell_6t_3 inst_cell_111_27 ( BL27, BLN27, WL111);
sram_cell_6t_3 inst_cell_111_26 ( BL26, BLN26, WL111);
sram_cell_6t_3 inst_cell_111_25 ( BL25, BLN25, WL111);
sram_cell_6t_3 inst_cell_111_24 ( BL24, BLN24, WL111);
sram_cell_6t_3 inst_cell_111_23 ( BL23, BLN23, WL111);
sram_cell_6t_3 inst_cell_111_22 ( BL22, BLN22, WL111);
sram_cell_6t_3 inst_cell_111_21 ( BL21, BLN21, WL111);
sram_cell_6t_3 inst_cell_111_20 ( BL20, BLN20, WL111);
sram_cell_6t_3 inst_cell_111_19 ( BL19, BLN19, WL111);
sram_cell_6t_3 inst_cell_111_18 ( BL18, BLN18, WL111);
sram_cell_6t_3 inst_cell_111_17 ( BL17, BLN17, WL111);
sram_cell_6t_3 inst_cell_111_16 ( BL16, BLN16, WL111);
sram_cell_6t_3 inst_cell_111_15 ( BL15, BLN15, WL111);
sram_cell_6t_3 inst_cell_111_14 ( BL14, BLN14, WL111);
sram_cell_6t_3 inst_cell_111_13 ( BL13, BLN13, WL111);
sram_cell_6t_3 inst_cell_111_12 ( BL12, BLN12, WL111);
sram_cell_6t_3 inst_cell_111_11 ( BL11, BLN11, WL111);
sram_cell_6t_3 inst_cell_111_10 ( BL10, BLN10, WL111);
sram_cell_6t_3 inst_cell_111_9 ( BL9, BLN9, WL111);
sram_cell_6t_3 inst_cell_111_8 ( BL8, BLN8, WL111);
sram_cell_6t_3 inst_cell_111_7 ( BL7, BLN7, WL111);
sram_cell_6t_3 inst_cell_111_6 ( BL6, BLN6, WL111);
sram_cell_6t_3 inst_cell_111_5 ( BL5, BLN5, WL111);
sram_cell_6t_3 inst_cell_111_4 ( BL4, BLN4, WL111);
sram_cell_6t_3 inst_cell_111_3 ( BL3, BLN3, WL111);
sram_cell_6t_3 inst_cell_111_2 ( BL2, BLN2, WL111);
sram_cell_6t_3 inst_cell_111_1 ( BL1, BLN1, WL111);
sram_cell_6t_3 inst_cell_111_0 ( BL0, BLN0, WL111);
sram_cell_6t_3 inst_cell_110_127 ( BL127, BLN127, WL110);
sram_cell_6t_3 inst_cell_110_126 ( BL126, BLN126, WL110);
sram_cell_6t_3 inst_cell_110_125 ( BL125, BLN125, WL110);
sram_cell_6t_3 inst_cell_110_124 ( BL124, BLN124, WL110);
sram_cell_6t_3 inst_cell_110_123 ( BL123, BLN123, WL110);
sram_cell_6t_3 inst_cell_110_122 ( BL122, BLN122, WL110);
sram_cell_6t_3 inst_cell_110_121 ( BL121, BLN121, WL110);
sram_cell_6t_3 inst_cell_110_120 ( BL120, BLN120, WL110);
sram_cell_6t_3 inst_cell_110_119 ( BL119, BLN119, WL110);
sram_cell_6t_3 inst_cell_110_118 ( BL118, BLN118, WL110);
sram_cell_6t_3 inst_cell_110_117 ( BL117, BLN117, WL110);
sram_cell_6t_3 inst_cell_110_116 ( BL116, BLN116, WL110);
sram_cell_6t_3 inst_cell_110_115 ( BL115, BLN115, WL110);
sram_cell_6t_3 inst_cell_110_114 ( BL114, BLN114, WL110);
sram_cell_6t_3 inst_cell_110_113 ( BL113, BLN113, WL110);
sram_cell_6t_3 inst_cell_110_112 ( BL112, BLN112, WL110);
sram_cell_6t_3 inst_cell_110_111 ( BL111, BLN111, WL110);
sram_cell_6t_3 inst_cell_110_110 ( BL110, BLN110, WL110);
sram_cell_6t_3 inst_cell_110_109 ( BL109, BLN109, WL110);
sram_cell_6t_3 inst_cell_110_108 ( BL108, BLN108, WL110);
sram_cell_6t_3 inst_cell_110_107 ( BL107, BLN107, WL110);
sram_cell_6t_3 inst_cell_110_106 ( BL106, BLN106, WL110);
sram_cell_6t_3 inst_cell_110_105 ( BL105, BLN105, WL110);
sram_cell_6t_3 inst_cell_110_104 ( BL104, BLN104, WL110);
sram_cell_6t_3 inst_cell_110_103 ( BL103, BLN103, WL110);
sram_cell_6t_3 inst_cell_110_102 ( BL102, BLN102, WL110);
sram_cell_6t_3 inst_cell_110_101 ( BL101, BLN101, WL110);
sram_cell_6t_3 inst_cell_110_100 ( BL100, BLN100, WL110);
sram_cell_6t_3 inst_cell_110_99 ( BL99, BLN99, WL110);
sram_cell_6t_3 inst_cell_110_98 ( BL98, BLN98, WL110);
sram_cell_6t_3 inst_cell_110_97 ( BL97, BLN97, WL110);
sram_cell_6t_3 inst_cell_110_96 ( BL96, BLN96, WL110);
sram_cell_6t_3 inst_cell_110_95 ( BL95, BLN95, WL110);
sram_cell_6t_3 inst_cell_110_94 ( BL94, BLN94, WL110);
sram_cell_6t_3 inst_cell_110_93 ( BL93, BLN93, WL110);
sram_cell_6t_3 inst_cell_110_92 ( BL92, BLN92, WL110);
sram_cell_6t_3 inst_cell_110_91 ( BL91, BLN91, WL110);
sram_cell_6t_3 inst_cell_110_90 ( BL90, BLN90, WL110);
sram_cell_6t_3 inst_cell_110_89 ( BL89, BLN89, WL110);
sram_cell_6t_3 inst_cell_110_88 ( BL88, BLN88, WL110);
sram_cell_6t_3 inst_cell_110_87 ( BL87, BLN87, WL110);
sram_cell_6t_3 inst_cell_110_86 ( BL86, BLN86, WL110);
sram_cell_6t_3 inst_cell_110_85 ( BL85, BLN85, WL110);
sram_cell_6t_3 inst_cell_110_84 ( BL84, BLN84, WL110);
sram_cell_6t_3 inst_cell_110_83 ( BL83, BLN83, WL110);
sram_cell_6t_3 inst_cell_110_82 ( BL82, BLN82, WL110);
sram_cell_6t_3 inst_cell_110_81 ( BL81, BLN81, WL110);
sram_cell_6t_3 inst_cell_110_80 ( BL80, BLN80, WL110);
sram_cell_6t_3 inst_cell_110_79 ( BL79, BLN79, WL110);
sram_cell_6t_3 inst_cell_110_78 ( BL78, BLN78, WL110);
sram_cell_6t_3 inst_cell_110_77 ( BL77, BLN77, WL110);
sram_cell_6t_3 inst_cell_110_76 ( BL76, BLN76, WL110);
sram_cell_6t_3 inst_cell_110_75 ( BL75, BLN75, WL110);
sram_cell_6t_3 inst_cell_110_74 ( BL74, BLN74, WL110);
sram_cell_6t_3 inst_cell_110_73 ( BL73, BLN73, WL110);
sram_cell_6t_3 inst_cell_110_72 ( BL72, BLN72, WL110);
sram_cell_6t_3 inst_cell_110_71 ( BL71, BLN71, WL110);
sram_cell_6t_3 inst_cell_110_70 ( BL70, BLN70, WL110);
sram_cell_6t_3 inst_cell_110_69 ( BL69, BLN69, WL110);
sram_cell_6t_3 inst_cell_110_68 ( BL68, BLN68, WL110);
sram_cell_6t_3 inst_cell_110_67 ( BL67, BLN67, WL110);
sram_cell_6t_3 inst_cell_110_66 ( BL66, BLN66, WL110);
sram_cell_6t_3 inst_cell_110_65 ( BL65, BLN65, WL110);
sram_cell_6t_3 inst_cell_110_64 ( BL64, BLN64, WL110);
sram_cell_6t_3 inst_cell_110_63 ( BL63, BLN63, WL110);
sram_cell_6t_3 inst_cell_110_62 ( BL62, BLN62, WL110);
sram_cell_6t_3 inst_cell_110_61 ( BL61, BLN61, WL110);
sram_cell_6t_3 inst_cell_110_60 ( BL60, BLN60, WL110);
sram_cell_6t_3 inst_cell_110_59 ( BL59, BLN59, WL110);
sram_cell_6t_3 inst_cell_110_58 ( BL58, BLN58, WL110);
sram_cell_6t_3 inst_cell_110_57 ( BL57, BLN57, WL110);
sram_cell_6t_3 inst_cell_110_56 ( BL56, BLN56, WL110);
sram_cell_6t_3 inst_cell_110_55 ( BL55, BLN55, WL110);
sram_cell_6t_3 inst_cell_110_54 ( BL54, BLN54, WL110);
sram_cell_6t_3 inst_cell_110_53 ( BL53, BLN53, WL110);
sram_cell_6t_3 inst_cell_110_52 ( BL52, BLN52, WL110);
sram_cell_6t_3 inst_cell_110_51 ( BL51, BLN51, WL110);
sram_cell_6t_3 inst_cell_110_50 ( BL50, BLN50, WL110);
sram_cell_6t_3 inst_cell_110_49 ( BL49, BLN49, WL110);
sram_cell_6t_3 inst_cell_110_48 ( BL48, BLN48, WL110);
sram_cell_6t_3 inst_cell_110_47 ( BL47, BLN47, WL110);
sram_cell_6t_3 inst_cell_110_46 ( BL46, BLN46, WL110);
sram_cell_6t_3 inst_cell_110_45 ( BL45, BLN45, WL110);
sram_cell_6t_3 inst_cell_110_44 ( BL44, BLN44, WL110);
sram_cell_6t_3 inst_cell_110_43 ( BL43, BLN43, WL110);
sram_cell_6t_3 inst_cell_110_42 ( BL42, BLN42, WL110);
sram_cell_6t_3 inst_cell_110_41 ( BL41, BLN41, WL110);
sram_cell_6t_3 inst_cell_110_40 ( BL40, BLN40, WL110);
sram_cell_6t_3 inst_cell_110_39 ( BL39, BLN39, WL110);
sram_cell_6t_3 inst_cell_110_38 ( BL38, BLN38, WL110);
sram_cell_6t_3 inst_cell_110_37 ( BL37, BLN37, WL110);
sram_cell_6t_3 inst_cell_110_36 ( BL36, BLN36, WL110);
sram_cell_6t_3 inst_cell_110_35 ( BL35, BLN35, WL110);
sram_cell_6t_3 inst_cell_110_34 ( BL34, BLN34, WL110);
sram_cell_6t_3 inst_cell_110_33 ( BL33, BLN33, WL110);
sram_cell_6t_3 inst_cell_110_32 ( BL32, BLN32, WL110);
sram_cell_6t_3 inst_cell_110_31 ( BL31, BLN31, WL110);
sram_cell_6t_3 inst_cell_110_30 ( BL30, BLN30, WL110);
sram_cell_6t_3 inst_cell_110_29 ( BL29, BLN29, WL110);
sram_cell_6t_3 inst_cell_110_28 ( BL28, BLN28, WL110);
sram_cell_6t_3 inst_cell_110_27 ( BL27, BLN27, WL110);
sram_cell_6t_3 inst_cell_110_26 ( BL26, BLN26, WL110);
sram_cell_6t_3 inst_cell_110_25 ( BL25, BLN25, WL110);
sram_cell_6t_3 inst_cell_110_24 ( BL24, BLN24, WL110);
sram_cell_6t_3 inst_cell_110_23 ( BL23, BLN23, WL110);
sram_cell_6t_3 inst_cell_110_22 ( BL22, BLN22, WL110);
sram_cell_6t_3 inst_cell_110_21 ( BL21, BLN21, WL110);
sram_cell_6t_3 inst_cell_110_20 ( BL20, BLN20, WL110);
sram_cell_6t_3 inst_cell_110_19 ( BL19, BLN19, WL110);
sram_cell_6t_3 inst_cell_110_18 ( BL18, BLN18, WL110);
sram_cell_6t_3 inst_cell_110_17 ( BL17, BLN17, WL110);
sram_cell_6t_3 inst_cell_110_16 ( BL16, BLN16, WL110);
sram_cell_6t_3 inst_cell_110_15 ( BL15, BLN15, WL110);
sram_cell_6t_3 inst_cell_110_14 ( BL14, BLN14, WL110);
sram_cell_6t_3 inst_cell_110_13 ( BL13, BLN13, WL110);
sram_cell_6t_3 inst_cell_110_12 ( BL12, BLN12, WL110);
sram_cell_6t_3 inst_cell_110_11 ( BL11, BLN11, WL110);
sram_cell_6t_3 inst_cell_110_10 ( BL10, BLN10, WL110);
sram_cell_6t_3 inst_cell_110_9 ( BL9, BLN9, WL110);
sram_cell_6t_3 inst_cell_110_8 ( BL8, BLN8, WL110);
sram_cell_6t_3 inst_cell_110_7 ( BL7, BLN7, WL110);
sram_cell_6t_3 inst_cell_110_6 ( BL6, BLN6, WL110);
sram_cell_6t_3 inst_cell_110_5 ( BL5, BLN5, WL110);
sram_cell_6t_3 inst_cell_110_4 ( BL4, BLN4, WL110);
sram_cell_6t_3 inst_cell_110_3 ( BL3, BLN3, WL110);
sram_cell_6t_3 inst_cell_110_2 ( BL2, BLN2, WL110);
sram_cell_6t_3 inst_cell_110_1 ( BL1, BLN1, WL110);
sram_cell_6t_3 inst_cell_110_0 ( BL0, BLN0, WL110);
sram_cell_6t_3 inst_cell_109_127 ( BL127, BLN127, WL109);
sram_cell_6t_3 inst_cell_109_126 ( BL126, BLN126, WL109);
sram_cell_6t_3 inst_cell_109_125 ( BL125, BLN125, WL109);
sram_cell_6t_3 inst_cell_109_124 ( BL124, BLN124, WL109);
sram_cell_6t_3 inst_cell_109_123 ( BL123, BLN123, WL109);
sram_cell_6t_3 inst_cell_109_122 ( BL122, BLN122, WL109);
sram_cell_6t_3 inst_cell_109_121 ( BL121, BLN121, WL109);
sram_cell_6t_3 inst_cell_109_120 ( BL120, BLN120, WL109);
sram_cell_6t_3 inst_cell_109_119 ( BL119, BLN119, WL109);
sram_cell_6t_3 inst_cell_109_118 ( BL118, BLN118, WL109);
sram_cell_6t_3 inst_cell_109_117 ( BL117, BLN117, WL109);
sram_cell_6t_3 inst_cell_109_116 ( BL116, BLN116, WL109);
sram_cell_6t_3 inst_cell_109_115 ( BL115, BLN115, WL109);
sram_cell_6t_3 inst_cell_109_114 ( BL114, BLN114, WL109);
sram_cell_6t_3 inst_cell_109_113 ( BL113, BLN113, WL109);
sram_cell_6t_3 inst_cell_109_112 ( BL112, BLN112, WL109);
sram_cell_6t_3 inst_cell_109_111 ( BL111, BLN111, WL109);
sram_cell_6t_3 inst_cell_109_110 ( BL110, BLN110, WL109);
sram_cell_6t_3 inst_cell_109_109 ( BL109, BLN109, WL109);
sram_cell_6t_3 inst_cell_109_108 ( BL108, BLN108, WL109);
sram_cell_6t_3 inst_cell_109_107 ( BL107, BLN107, WL109);
sram_cell_6t_3 inst_cell_109_106 ( BL106, BLN106, WL109);
sram_cell_6t_3 inst_cell_109_105 ( BL105, BLN105, WL109);
sram_cell_6t_3 inst_cell_109_104 ( BL104, BLN104, WL109);
sram_cell_6t_3 inst_cell_109_103 ( BL103, BLN103, WL109);
sram_cell_6t_3 inst_cell_109_102 ( BL102, BLN102, WL109);
sram_cell_6t_3 inst_cell_109_101 ( BL101, BLN101, WL109);
sram_cell_6t_3 inst_cell_109_100 ( BL100, BLN100, WL109);
sram_cell_6t_3 inst_cell_109_99 ( BL99, BLN99, WL109);
sram_cell_6t_3 inst_cell_109_98 ( BL98, BLN98, WL109);
sram_cell_6t_3 inst_cell_109_97 ( BL97, BLN97, WL109);
sram_cell_6t_3 inst_cell_109_96 ( BL96, BLN96, WL109);
sram_cell_6t_3 inst_cell_109_95 ( BL95, BLN95, WL109);
sram_cell_6t_3 inst_cell_109_94 ( BL94, BLN94, WL109);
sram_cell_6t_3 inst_cell_109_93 ( BL93, BLN93, WL109);
sram_cell_6t_3 inst_cell_109_92 ( BL92, BLN92, WL109);
sram_cell_6t_3 inst_cell_109_91 ( BL91, BLN91, WL109);
sram_cell_6t_3 inst_cell_109_90 ( BL90, BLN90, WL109);
sram_cell_6t_3 inst_cell_109_89 ( BL89, BLN89, WL109);
sram_cell_6t_3 inst_cell_109_88 ( BL88, BLN88, WL109);
sram_cell_6t_3 inst_cell_109_87 ( BL87, BLN87, WL109);
sram_cell_6t_3 inst_cell_109_86 ( BL86, BLN86, WL109);
sram_cell_6t_3 inst_cell_109_85 ( BL85, BLN85, WL109);
sram_cell_6t_3 inst_cell_109_84 ( BL84, BLN84, WL109);
sram_cell_6t_3 inst_cell_109_83 ( BL83, BLN83, WL109);
sram_cell_6t_3 inst_cell_109_82 ( BL82, BLN82, WL109);
sram_cell_6t_3 inst_cell_109_81 ( BL81, BLN81, WL109);
sram_cell_6t_3 inst_cell_109_80 ( BL80, BLN80, WL109);
sram_cell_6t_3 inst_cell_109_79 ( BL79, BLN79, WL109);
sram_cell_6t_3 inst_cell_109_78 ( BL78, BLN78, WL109);
sram_cell_6t_3 inst_cell_109_77 ( BL77, BLN77, WL109);
sram_cell_6t_3 inst_cell_109_76 ( BL76, BLN76, WL109);
sram_cell_6t_3 inst_cell_109_75 ( BL75, BLN75, WL109);
sram_cell_6t_3 inst_cell_109_74 ( BL74, BLN74, WL109);
sram_cell_6t_3 inst_cell_109_73 ( BL73, BLN73, WL109);
sram_cell_6t_3 inst_cell_109_72 ( BL72, BLN72, WL109);
sram_cell_6t_3 inst_cell_109_71 ( BL71, BLN71, WL109);
sram_cell_6t_3 inst_cell_109_70 ( BL70, BLN70, WL109);
sram_cell_6t_3 inst_cell_109_69 ( BL69, BLN69, WL109);
sram_cell_6t_3 inst_cell_109_68 ( BL68, BLN68, WL109);
sram_cell_6t_3 inst_cell_109_67 ( BL67, BLN67, WL109);
sram_cell_6t_3 inst_cell_109_66 ( BL66, BLN66, WL109);
sram_cell_6t_3 inst_cell_109_65 ( BL65, BLN65, WL109);
sram_cell_6t_3 inst_cell_109_64 ( BL64, BLN64, WL109);
sram_cell_6t_3 inst_cell_109_63 ( BL63, BLN63, WL109);
sram_cell_6t_3 inst_cell_109_62 ( BL62, BLN62, WL109);
sram_cell_6t_3 inst_cell_109_61 ( BL61, BLN61, WL109);
sram_cell_6t_3 inst_cell_109_60 ( BL60, BLN60, WL109);
sram_cell_6t_3 inst_cell_109_59 ( BL59, BLN59, WL109);
sram_cell_6t_3 inst_cell_109_58 ( BL58, BLN58, WL109);
sram_cell_6t_3 inst_cell_109_57 ( BL57, BLN57, WL109);
sram_cell_6t_3 inst_cell_109_56 ( BL56, BLN56, WL109);
sram_cell_6t_3 inst_cell_109_55 ( BL55, BLN55, WL109);
sram_cell_6t_3 inst_cell_109_54 ( BL54, BLN54, WL109);
sram_cell_6t_3 inst_cell_109_53 ( BL53, BLN53, WL109);
sram_cell_6t_3 inst_cell_109_52 ( BL52, BLN52, WL109);
sram_cell_6t_3 inst_cell_109_51 ( BL51, BLN51, WL109);
sram_cell_6t_3 inst_cell_109_50 ( BL50, BLN50, WL109);
sram_cell_6t_3 inst_cell_109_49 ( BL49, BLN49, WL109);
sram_cell_6t_3 inst_cell_109_48 ( BL48, BLN48, WL109);
sram_cell_6t_3 inst_cell_109_47 ( BL47, BLN47, WL109);
sram_cell_6t_3 inst_cell_109_46 ( BL46, BLN46, WL109);
sram_cell_6t_3 inst_cell_109_45 ( BL45, BLN45, WL109);
sram_cell_6t_3 inst_cell_109_44 ( BL44, BLN44, WL109);
sram_cell_6t_3 inst_cell_109_43 ( BL43, BLN43, WL109);
sram_cell_6t_3 inst_cell_109_42 ( BL42, BLN42, WL109);
sram_cell_6t_3 inst_cell_109_41 ( BL41, BLN41, WL109);
sram_cell_6t_3 inst_cell_109_40 ( BL40, BLN40, WL109);
sram_cell_6t_3 inst_cell_109_39 ( BL39, BLN39, WL109);
sram_cell_6t_3 inst_cell_109_38 ( BL38, BLN38, WL109);
sram_cell_6t_3 inst_cell_109_37 ( BL37, BLN37, WL109);
sram_cell_6t_3 inst_cell_109_36 ( BL36, BLN36, WL109);
sram_cell_6t_3 inst_cell_109_35 ( BL35, BLN35, WL109);
sram_cell_6t_3 inst_cell_109_34 ( BL34, BLN34, WL109);
sram_cell_6t_3 inst_cell_109_33 ( BL33, BLN33, WL109);
sram_cell_6t_3 inst_cell_109_32 ( BL32, BLN32, WL109);
sram_cell_6t_3 inst_cell_109_31 ( BL31, BLN31, WL109);
sram_cell_6t_3 inst_cell_109_30 ( BL30, BLN30, WL109);
sram_cell_6t_3 inst_cell_109_29 ( BL29, BLN29, WL109);
sram_cell_6t_3 inst_cell_109_28 ( BL28, BLN28, WL109);
sram_cell_6t_3 inst_cell_109_27 ( BL27, BLN27, WL109);
sram_cell_6t_3 inst_cell_109_26 ( BL26, BLN26, WL109);
sram_cell_6t_3 inst_cell_109_25 ( BL25, BLN25, WL109);
sram_cell_6t_3 inst_cell_109_24 ( BL24, BLN24, WL109);
sram_cell_6t_3 inst_cell_109_23 ( BL23, BLN23, WL109);
sram_cell_6t_3 inst_cell_109_22 ( BL22, BLN22, WL109);
sram_cell_6t_3 inst_cell_109_21 ( BL21, BLN21, WL109);
sram_cell_6t_3 inst_cell_109_20 ( BL20, BLN20, WL109);
sram_cell_6t_3 inst_cell_109_19 ( BL19, BLN19, WL109);
sram_cell_6t_3 inst_cell_109_18 ( BL18, BLN18, WL109);
sram_cell_6t_3 inst_cell_109_17 ( BL17, BLN17, WL109);
sram_cell_6t_3 inst_cell_109_16 ( BL16, BLN16, WL109);
sram_cell_6t_3 inst_cell_109_15 ( BL15, BLN15, WL109);
sram_cell_6t_3 inst_cell_109_14 ( BL14, BLN14, WL109);
sram_cell_6t_3 inst_cell_109_13 ( BL13, BLN13, WL109);
sram_cell_6t_3 inst_cell_109_12 ( BL12, BLN12, WL109);
sram_cell_6t_3 inst_cell_109_11 ( BL11, BLN11, WL109);
sram_cell_6t_3 inst_cell_109_10 ( BL10, BLN10, WL109);
sram_cell_6t_3 inst_cell_109_9 ( BL9, BLN9, WL109);
sram_cell_6t_3 inst_cell_109_8 ( BL8, BLN8, WL109);
sram_cell_6t_3 inst_cell_109_7 ( BL7, BLN7, WL109);
sram_cell_6t_3 inst_cell_109_6 ( BL6, BLN6, WL109);
sram_cell_6t_3 inst_cell_109_5 ( BL5, BLN5, WL109);
sram_cell_6t_3 inst_cell_109_4 ( BL4, BLN4, WL109);
sram_cell_6t_3 inst_cell_109_3 ( BL3, BLN3, WL109);
sram_cell_6t_3 inst_cell_109_2 ( BL2, BLN2, WL109);
sram_cell_6t_3 inst_cell_109_1 ( BL1, BLN1, WL109);
sram_cell_6t_3 inst_cell_109_0 ( BL0, BLN0, WL109);
sram_cell_6t_3 inst_cell_108_127 ( BL127, BLN127, WL108);
sram_cell_6t_3 inst_cell_108_126 ( BL126, BLN126, WL108);
sram_cell_6t_3 inst_cell_108_125 ( BL125, BLN125, WL108);
sram_cell_6t_3 inst_cell_108_124 ( BL124, BLN124, WL108);
sram_cell_6t_3 inst_cell_108_123 ( BL123, BLN123, WL108);
sram_cell_6t_3 inst_cell_108_122 ( BL122, BLN122, WL108);
sram_cell_6t_3 inst_cell_108_121 ( BL121, BLN121, WL108);
sram_cell_6t_3 inst_cell_108_120 ( BL120, BLN120, WL108);
sram_cell_6t_3 inst_cell_108_119 ( BL119, BLN119, WL108);
sram_cell_6t_3 inst_cell_108_118 ( BL118, BLN118, WL108);
sram_cell_6t_3 inst_cell_108_117 ( BL117, BLN117, WL108);
sram_cell_6t_3 inst_cell_108_116 ( BL116, BLN116, WL108);
sram_cell_6t_3 inst_cell_108_115 ( BL115, BLN115, WL108);
sram_cell_6t_3 inst_cell_108_114 ( BL114, BLN114, WL108);
sram_cell_6t_3 inst_cell_108_113 ( BL113, BLN113, WL108);
sram_cell_6t_3 inst_cell_108_112 ( BL112, BLN112, WL108);
sram_cell_6t_3 inst_cell_108_111 ( BL111, BLN111, WL108);
sram_cell_6t_3 inst_cell_108_110 ( BL110, BLN110, WL108);
sram_cell_6t_3 inst_cell_108_109 ( BL109, BLN109, WL108);
sram_cell_6t_3 inst_cell_108_108 ( BL108, BLN108, WL108);
sram_cell_6t_3 inst_cell_108_107 ( BL107, BLN107, WL108);
sram_cell_6t_3 inst_cell_108_106 ( BL106, BLN106, WL108);
sram_cell_6t_3 inst_cell_108_105 ( BL105, BLN105, WL108);
sram_cell_6t_3 inst_cell_108_104 ( BL104, BLN104, WL108);
sram_cell_6t_3 inst_cell_108_103 ( BL103, BLN103, WL108);
sram_cell_6t_3 inst_cell_108_102 ( BL102, BLN102, WL108);
sram_cell_6t_3 inst_cell_108_101 ( BL101, BLN101, WL108);
sram_cell_6t_3 inst_cell_108_100 ( BL100, BLN100, WL108);
sram_cell_6t_3 inst_cell_108_99 ( BL99, BLN99, WL108);
sram_cell_6t_3 inst_cell_108_98 ( BL98, BLN98, WL108);
sram_cell_6t_3 inst_cell_108_97 ( BL97, BLN97, WL108);
sram_cell_6t_3 inst_cell_108_96 ( BL96, BLN96, WL108);
sram_cell_6t_3 inst_cell_108_95 ( BL95, BLN95, WL108);
sram_cell_6t_3 inst_cell_108_94 ( BL94, BLN94, WL108);
sram_cell_6t_3 inst_cell_108_93 ( BL93, BLN93, WL108);
sram_cell_6t_3 inst_cell_108_92 ( BL92, BLN92, WL108);
sram_cell_6t_3 inst_cell_108_91 ( BL91, BLN91, WL108);
sram_cell_6t_3 inst_cell_108_90 ( BL90, BLN90, WL108);
sram_cell_6t_3 inst_cell_108_89 ( BL89, BLN89, WL108);
sram_cell_6t_3 inst_cell_108_88 ( BL88, BLN88, WL108);
sram_cell_6t_3 inst_cell_108_87 ( BL87, BLN87, WL108);
sram_cell_6t_3 inst_cell_108_86 ( BL86, BLN86, WL108);
sram_cell_6t_3 inst_cell_108_85 ( BL85, BLN85, WL108);
sram_cell_6t_3 inst_cell_108_84 ( BL84, BLN84, WL108);
sram_cell_6t_3 inst_cell_108_83 ( BL83, BLN83, WL108);
sram_cell_6t_3 inst_cell_108_82 ( BL82, BLN82, WL108);
sram_cell_6t_3 inst_cell_108_81 ( BL81, BLN81, WL108);
sram_cell_6t_3 inst_cell_108_80 ( BL80, BLN80, WL108);
sram_cell_6t_3 inst_cell_108_79 ( BL79, BLN79, WL108);
sram_cell_6t_3 inst_cell_108_78 ( BL78, BLN78, WL108);
sram_cell_6t_3 inst_cell_108_77 ( BL77, BLN77, WL108);
sram_cell_6t_3 inst_cell_108_76 ( BL76, BLN76, WL108);
sram_cell_6t_3 inst_cell_108_75 ( BL75, BLN75, WL108);
sram_cell_6t_3 inst_cell_108_74 ( BL74, BLN74, WL108);
sram_cell_6t_3 inst_cell_108_73 ( BL73, BLN73, WL108);
sram_cell_6t_3 inst_cell_108_72 ( BL72, BLN72, WL108);
sram_cell_6t_3 inst_cell_108_71 ( BL71, BLN71, WL108);
sram_cell_6t_3 inst_cell_108_70 ( BL70, BLN70, WL108);
sram_cell_6t_3 inst_cell_108_69 ( BL69, BLN69, WL108);
sram_cell_6t_3 inst_cell_108_68 ( BL68, BLN68, WL108);
sram_cell_6t_3 inst_cell_108_67 ( BL67, BLN67, WL108);
sram_cell_6t_3 inst_cell_108_66 ( BL66, BLN66, WL108);
sram_cell_6t_3 inst_cell_108_65 ( BL65, BLN65, WL108);
sram_cell_6t_3 inst_cell_108_64 ( BL64, BLN64, WL108);
sram_cell_6t_3 inst_cell_108_63 ( BL63, BLN63, WL108);
sram_cell_6t_3 inst_cell_108_62 ( BL62, BLN62, WL108);
sram_cell_6t_3 inst_cell_108_61 ( BL61, BLN61, WL108);
sram_cell_6t_3 inst_cell_108_60 ( BL60, BLN60, WL108);
sram_cell_6t_3 inst_cell_108_59 ( BL59, BLN59, WL108);
sram_cell_6t_3 inst_cell_108_58 ( BL58, BLN58, WL108);
sram_cell_6t_3 inst_cell_108_57 ( BL57, BLN57, WL108);
sram_cell_6t_3 inst_cell_108_56 ( BL56, BLN56, WL108);
sram_cell_6t_3 inst_cell_108_55 ( BL55, BLN55, WL108);
sram_cell_6t_3 inst_cell_108_54 ( BL54, BLN54, WL108);
sram_cell_6t_3 inst_cell_108_53 ( BL53, BLN53, WL108);
sram_cell_6t_3 inst_cell_108_52 ( BL52, BLN52, WL108);
sram_cell_6t_3 inst_cell_108_51 ( BL51, BLN51, WL108);
sram_cell_6t_3 inst_cell_108_50 ( BL50, BLN50, WL108);
sram_cell_6t_3 inst_cell_108_49 ( BL49, BLN49, WL108);
sram_cell_6t_3 inst_cell_108_48 ( BL48, BLN48, WL108);
sram_cell_6t_3 inst_cell_108_47 ( BL47, BLN47, WL108);
sram_cell_6t_3 inst_cell_108_46 ( BL46, BLN46, WL108);
sram_cell_6t_3 inst_cell_108_45 ( BL45, BLN45, WL108);
sram_cell_6t_3 inst_cell_108_44 ( BL44, BLN44, WL108);
sram_cell_6t_3 inst_cell_108_43 ( BL43, BLN43, WL108);
sram_cell_6t_3 inst_cell_108_42 ( BL42, BLN42, WL108);
sram_cell_6t_3 inst_cell_108_41 ( BL41, BLN41, WL108);
sram_cell_6t_3 inst_cell_108_40 ( BL40, BLN40, WL108);
sram_cell_6t_3 inst_cell_108_39 ( BL39, BLN39, WL108);
sram_cell_6t_3 inst_cell_108_38 ( BL38, BLN38, WL108);
sram_cell_6t_3 inst_cell_108_37 ( BL37, BLN37, WL108);
sram_cell_6t_3 inst_cell_108_36 ( BL36, BLN36, WL108);
sram_cell_6t_3 inst_cell_108_35 ( BL35, BLN35, WL108);
sram_cell_6t_3 inst_cell_108_34 ( BL34, BLN34, WL108);
sram_cell_6t_3 inst_cell_108_33 ( BL33, BLN33, WL108);
sram_cell_6t_3 inst_cell_108_32 ( BL32, BLN32, WL108);
sram_cell_6t_3 inst_cell_108_31 ( BL31, BLN31, WL108);
sram_cell_6t_3 inst_cell_108_30 ( BL30, BLN30, WL108);
sram_cell_6t_3 inst_cell_108_29 ( BL29, BLN29, WL108);
sram_cell_6t_3 inst_cell_108_28 ( BL28, BLN28, WL108);
sram_cell_6t_3 inst_cell_108_27 ( BL27, BLN27, WL108);
sram_cell_6t_3 inst_cell_108_26 ( BL26, BLN26, WL108);
sram_cell_6t_3 inst_cell_108_25 ( BL25, BLN25, WL108);
sram_cell_6t_3 inst_cell_108_24 ( BL24, BLN24, WL108);
sram_cell_6t_3 inst_cell_108_23 ( BL23, BLN23, WL108);
sram_cell_6t_3 inst_cell_108_22 ( BL22, BLN22, WL108);
sram_cell_6t_3 inst_cell_108_21 ( BL21, BLN21, WL108);
sram_cell_6t_3 inst_cell_108_20 ( BL20, BLN20, WL108);
sram_cell_6t_3 inst_cell_108_19 ( BL19, BLN19, WL108);
sram_cell_6t_3 inst_cell_108_18 ( BL18, BLN18, WL108);
sram_cell_6t_3 inst_cell_108_17 ( BL17, BLN17, WL108);
sram_cell_6t_3 inst_cell_108_16 ( BL16, BLN16, WL108);
sram_cell_6t_3 inst_cell_108_15 ( BL15, BLN15, WL108);
sram_cell_6t_3 inst_cell_108_14 ( BL14, BLN14, WL108);
sram_cell_6t_3 inst_cell_108_13 ( BL13, BLN13, WL108);
sram_cell_6t_3 inst_cell_108_12 ( BL12, BLN12, WL108);
sram_cell_6t_3 inst_cell_108_11 ( BL11, BLN11, WL108);
sram_cell_6t_3 inst_cell_108_10 ( BL10, BLN10, WL108);
sram_cell_6t_3 inst_cell_108_9 ( BL9, BLN9, WL108);
sram_cell_6t_3 inst_cell_108_8 ( BL8, BLN8, WL108);
sram_cell_6t_3 inst_cell_108_7 ( BL7, BLN7, WL108);
sram_cell_6t_3 inst_cell_108_6 ( BL6, BLN6, WL108);
sram_cell_6t_3 inst_cell_108_5 ( BL5, BLN5, WL108);
sram_cell_6t_3 inst_cell_108_4 ( BL4, BLN4, WL108);
sram_cell_6t_3 inst_cell_108_3 ( BL3, BLN3, WL108);
sram_cell_6t_3 inst_cell_108_2 ( BL2, BLN2, WL108);
sram_cell_6t_3 inst_cell_108_1 ( BL1, BLN1, WL108);
sram_cell_6t_3 inst_cell_108_0 ( BL0, BLN0, WL108);
sram_cell_6t_3 inst_cell_107_127 ( BL127, BLN127, WL107);
sram_cell_6t_3 inst_cell_107_126 ( BL126, BLN126, WL107);
sram_cell_6t_3 inst_cell_107_125 ( BL125, BLN125, WL107);
sram_cell_6t_3 inst_cell_107_124 ( BL124, BLN124, WL107);
sram_cell_6t_3 inst_cell_107_123 ( BL123, BLN123, WL107);
sram_cell_6t_3 inst_cell_107_122 ( BL122, BLN122, WL107);
sram_cell_6t_3 inst_cell_107_121 ( BL121, BLN121, WL107);
sram_cell_6t_3 inst_cell_107_120 ( BL120, BLN120, WL107);
sram_cell_6t_3 inst_cell_107_119 ( BL119, BLN119, WL107);
sram_cell_6t_3 inst_cell_107_118 ( BL118, BLN118, WL107);
sram_cell_6t_3 inst_cell_107_117 ( BL117, BLN117, WL107);
sram_cell_6t_3 inst_cell_107_116 ( BL116, BLN116, WL107);
sram_cell_6t_3 inst_cell_107_115 ( BL115, BLN115, WL107);
sram_cell_6t_3 inst_cell_107_114 ( BL114, BLN114, WL107);
sram_cell_6t_3 inst_cell_107_113 ( BL113, BLN113, WL107);
sram_cell_6t_3 inst_cell_107_112 ( BL112, BLN112, WL107);
sram_cell_6t_3 inst_cell_107_111 ( BL111, BLN111, WL107);
sram_cell_6t_3 inst_cell_107_110 ( BL110, BLN110, WL107);
sram_cell_6t_3 inst_cell_107_109 ( BL109, BLN109, WL107);
sram_cell_6t_3 inst_cell_107_108 ( BL108, BLN108, WL107);
sram_cell_6t_3 inst_cell_107_107 ( BL107, BLN107, WL107);
sram_cell_6t_3 inst_cell_107_106 ( BL106, BLN106, WL107);
sram_cell_6t_3 inst_cell_107_105 ( BL105, BLN105, WL107);
sram_cell_6t_3 inst_cell_107_104 ( BL104, BLN104, WL107);
sram_cell_6t_3 inst_cell_107_103 ( BL103, BLN103, WL107);
sram_cell_6t_3 inst_cell_107_102 ( BL102, BLN102, WL107);
sram_cell_6t_3 inst_cell_107_101 ( BL101, BLN101, WL107);
sram_cell_6t_3 inst_cell_107_100 ( BL100, BLN100, WL107);
sram_cell_6t_3 inst_cell_107_99 ( BL99, BLN99, WL107);
sram_cell_6t_3 inst_cell_107_98 ( BL98, BLN98, WL107);
sram_cell_6t_3 inst_cell_107_97 ( BL97, BLN97, WL107);
sram_cell_6t_3 inst_cell_107_96 ( BL96, BLN96, WL107);
sram_cell_6t_3 inst_cell_107_95 ( BL95, BLN95, WL107);
sram_cell_6t_3 inst_cell_107_94 ( BL94, BLN94, WL107);
sram_cell_6t_3 inst_cell_107_93 ( BL93, BLN93, WL107);
sram_cell_6t_3 inst_cell_107_92 ( BL92, BLN92, WL107);
sram_cell_6t_3 inst_cell_107_91 ( BL91, BLN91, WL107);
sram_cell_6t_3 inst_cell_107_90 ( BL90, BLN90, WL107);
sram_cell_6t_3 inst_cell_107_89 ( BL89, BLN89, WL107);
sram_cell_6t_3 inst_cell_107_88 ( BL88, BLN88, WL107);
sram_cell_6t_3 inst_cell_107_87 ( BL87, BLN87, WL107);
sram_cell_6t_3 inst_cell_107_86 ( BL86, BLN86, WL107);
sram_cell_6t_3 inst_cell_107_85 ( BL85, BLN85, WL107);
sram_cell_6t_3 inst_cell_107_84 ( BL84, BLN84, WL107);
sram_cell_6t_3 inst_cell_107_83 ( BL83, BLN83, WL107);
sram_cell_6t_3 inst_cell_107_82 ( BL82, BLN82, WL107);
sram_cell_6t_3 inst_cell_107_81 ( BL81, BLN81, WL107);
sram_cell_6t_3 inst_cell_107_80 ( BL80, BLN80, WL107);
sram_cell_6t_3 inst_cell_107_79 ( BL79, BLN79, WL107);
sram_cell_6t_3 inst_cell_107_78 ( BL78, BLN78, WL107);
sram_cell_6t_3 inst_cell_107_77 ( BL77, BLN77, WL107);
sram_cell_6t_3 inst_cell_107_76 ( BL76, BLN76, WL107);
sram_cell_6t_3 inst_cell_107_75 ( BL75, BLN75, WL107);
sram_cell_6t_3 inst_cell_107_74 ( BL74, BLN74, WL107);
sram_cell_6t_3 inst_cell_107_73 ( BL73, BLN73, WL107);
sram_cell_6t_3 inst_cell_107_72 ( BL72, BLN72, WL107);
sram_cell_6t_3 inst_cell_107_71 ( BL71, BLN71, WL107);
sram_cell_6t_3 inst_cell_107_70 ( BL70, BLN70, WL107);
sram_cell_6t_3 inst_cell_107_69 ( BL69, BLN69, WL107);
sram_cell_6t_3 inst_cell_107_68 ( BL68, BLN68, WL107);
sram_cell_6t_3 inst_cell_107_67 ( BL67, BLN67, WL107);
sram_cell_6t_3 inst_cell_107_66 ( BL66, BLN66, WL107);
sram_cell_6t_3 inst_cell_107_65 ( BL65, BLN65, WL107);
sram_cell_6t_3 inst_cell_107_64 ( BL64, BLN64, WL107);
sram_cell_6t_3 inst_cell_107_63 ( BL63, BLN63, WL107);
sram_cell_6t_3 inst_cell_107_62 ( BL62, BLN62, WL107);
sram_cell_6t_3 inst_cell_107_61 ( BL61, BLN61, WL107);
sram_cell_6t_3 inst_cell_107_60 ( BL60, BLN60, WL107);
sram_cell_6t_3 inst_cell_107_59 ( BL59, BLN59, WL107);
sram_cell_6t_3 inst_cell_107_58 ( BL58, BLN58, WL107);
sram_cell_6t_3 inst_cell_107_57 ( BL57, BLN57, WL107);
sram_cell_6t_3 inst_cell_107_56 ( BL56, BLN56, WL107);
sram_cell_6t_3 inst_cell_107_55 ( BL55, BLN55, WL107);
sram_cell_6t_3 inst_cell_107_54 ( BL54, BLN54, WL107);
sram_cell_6t_3 inst_cell_107_53 ( BL53, BLN53, WL107);
sram_cell_6t_3 inst_cell_107_52 ( BL52, BLN52, WL107);
sram_cell_6t_3 inst_cell_107_51 ( BL51, BLN51, WL107);
sram_cell_6t_3 inst_cell_107_50 ( BL50, BLN50, WL107);
sram_cell_6t_3 inst_cell_107_49 ( BL49, BLN49, WL107);
sram_cell_6t_3 inst_cell_107_48 ( BL48, BLN48, WL107);
sram_cell_6t_3 inst_cell_107_47 ( BL47, BLN47, WL107);
sram_cell_6t_3 inst_cell_107_46 ( BL46, BLN46, WL107);
sram_cell_6t_3 inst_cell_107_45 ( BL45, BLN45, WL107);
sram_cell_6t_3 inst_cell_107_44 ( BL44, BLN44, WL107);
sram_cell_6t_3 inst_cell_107_43 ( BL43, BLN43, WL107);
sram_cell_6t_3 inst_cell_107_42 ( BL42, BLN42, WL107);
sram_cell_6t_3 inst_cell_107_41 ( BL41, BLN41, WL107);
sram_cell_6t_3 inst_cell_107_40 ( BL40, BLN40, WL107);
sram_cell_6t_3 inst_cell_107_39 ( BL39, BLN39, WL107);
sram_cell_6t_3 inst_cell_107_38 ( BL38, BLN38, WL107);
sram_cell_6t_3 inst_cell_107_37 ( BL37, BLN37, WL107);
sram_cell_6t_3 inst_cell_107_36 ( BL36, BLN36, WL107);
sram_cell_6t_3 inst_cell_107_35 ( BL35, BLN35, WL107);
sram_cell_6t_3 inst_cell_107_34 ( BL34, BLN34, WL107);
sram_cell_6t_3 inst_cell_107_33 ( BL33, BLN33, WL107);
sram_cell_6t_3 inst_cell_107_32 ( BL32, BLN32, WL107);
sram_cell_6t_3 inst_cell_107_31 ( BL31, BLN31, WL107);
sram_cell_6t_3 inst_cell_107_30 ( BL30, BLN30, WL107);
sram_cell_6t_3 inst_cell_107_29 ( BL29, BLN29, WL107);
sram_cell_6t_3 inst_cell_107_28 ( BL28, BLN28, WL107);
sram_cell_6t_3 inst_cell_107_27 ( BL27, BLN27, WL107);
sram_cell_6t_3 inst_cell_107_26 ( BL26, BLN26, WL107);
sram_cell_6t_3 inst_cell_107_25 ( BL25, BLN25, WL107);
sram_cell_6t_3 inst_cell_107_24 ( BL24, BLN24, WL107);
sram_cell_6t_3 inst_cell_107_23 ( BL23, BLN23, WL107);
sram_cell_6t_3 inst_cell_107_22 ( BL22, BLN22, WL107);
sram_cell_6t_3 inst_cell_107_21 ( BL21, BLN21, WL107);
sram_cell_6t_3 inst_cell_107_20 ( BL20, BLN20, WL107);
sram_cell_6t_3 inst_cell_107_19 ( BL19, BLN19, WL107);
sram_cell_6t_3 inst_cell_107_18 ( BL18, BLN18, WL107);
sram_cell_6t_3 inst_cell_107_17 ( BL17, BLN17, WL107);
sram_cell_6t_3 inst_cell_107_16 ( BL16, BLN16, WL107);
sram_cell_6t_3 inst_cell_107_15 ( BL15, BLN15, WL107);
sram_cell_6t_3 inst_cell_107_14 ( BL14, BLN14, WL107);
sram_cell_6t_3 inst_cell_107_13 ( BL13, BLN13, WL107);
sram_cell_6t_3 inst_cell_107_12 ( BL12, BLN12, WL107);
sram_cell_6t_3 inst_cell_107_11 ( BL11, BLN11, WL107);
sram_cell_6t_3 inst_cell_107_10 ( BL10, BLN10, WL107);
sram_cell_6t_3 inst_cell_107_9 ( BL9, BLN9, WL107);
sram_cell_6t_3 inst_cell_107_8 ( BL8, BLN8, WL107);
sram_cell_6t_3 inst_cell_107_7 ( BL7, BLN7, WL107);
sram_cell_6t_3 inst_cell_107_6 ( BL6, BLN6, WL107);
sram_cell_6t_3 inst_cell_107_5 ( BL5, BLN5, WL107);
sram_cell_6t_3 inst_cell_107_4 ( BL4, BLN4, WL107);
sram_cell_6t_3 inst_cell_107_3 ( BL3, BLN3, WL107);
sram_cell_6t_3 inst_cell_107_2 ( BL2, BLN2, WL107);
sram_cell_6t_3 inst_cell_107_1 ( BL1, BLN1, WL107);
sram_cell_6t_3 inst_cell_107_0 ( BL0, BLN0, WL107);
sram_cell_6t_3 inst_cell_106_127 ( BL127, BLN127, WL106);
sram_cell_6t_3 inst_cell_106_126 ( BL126, BLN126, WL106);
sram_cell_6t_3 inst_cell_106_125 ( BL125, BLN125, WL106);
sram_cell_6t_3 inst_cell_106_124 ( BL124, BLN124, WL106);
sram_cell_6t_3 inst_cell_106_123 ( BL123, BLN123, WL106);
sram_cell_6t_3 inst_cell_106_122 ( BL122, BLN122, WL106);
sram_cell_6t_3 inst_cell_106_121 ( BL121, BLN121, WL106);
sram_cell_6t_3 inst_cell_106_120 ( BL120, BLN120, WL106);
sram_cell_6t_3 inst_cell_106_119 ( BL119, BLN119, WL106);
sram_cell_6t_3 inst_cell_106_118 ( BL118, BLN118, WL106);
sram_cell_6t_3 inst_cell_106_117 ( BL117, BLN117, WL106);
sram_cell_6t_3 inst_cell_106_116 ( BL116, BLN116, WL106);
sram_cell_6t_3 inst_cell_106_115 ( BL115, BLN115, WL106);
sram_cell_6t_3 inst_cell_106_114 ( BL114, BLN114, WL106);
sram_cell_6t_3 inst_cell_106_113 ( BL113, BLN113, WL106);
sram_cell_6t_3 inst_cell_106_112 ( BL112, BLN112, WL106);
sram_cell_6t_3 inst_cell_106_111 ( BL111, BLN111, WL106);
sram_cell_6t_3 inst_cell_106_110 ( BL110, BLN110, WL106);
sram_cell_6t_3 inst_cell_106_109 ( BL109, BLN109, WL106);
sram_cell_6t_3 inst_cell_106_108 ( BL108, BLN108, WL106);
sram_cell_6t_3 inst_cell_106_107 ( BL107, BLN107, WL106);
sram_cell_6t_3 inst_cell_106_106 ( BL106, BLN106, WL106);
sram_cell_6t_3 inst_cell_106_105 ( BL105, BLN105, WL106);
sram_cell_6t_3 inst_cell_106_104 ( BL104, BLN104, WL106);
sram_cell_6t_3 inst_cell_106_103 ( BL103, BLN103, WL106);
sram_cell_6t_3 inst_cell_106_102 ( BL102, BLN102, WL106);
sram_cell_6t_3 inst_cell_106_101 ( BL101, BLN101, WL106);
sram_cell_6t_3 inst_cell_106_100 ( BL100, BLN100, WL106);
sram_cell_6t_3 inst_cell_106_99 ( BL99, BLN99, WL106);
sram_cell_6t_3 inst_cell_106_98 ( BL98, BLN98, WL106);
sram_cell_6t_3 inst_cell_106_97 ( BL97, BLN97, WL106);
sram_cell_6t_3 inst_cell_106_96 ( BL96, BLN96, WL106);
sram_cell_6t_3 inst_cell_106_95 ( BL95, BLN95, WL106);
sram_cell_6t_3 inst_cell_106_94 ( BL94, BLN94, WL106);
sram_cell_6t_3 inst_cell_106_93 ( BL93, BLN93, WL106);
sram_cell_6t_3 inst_cell_106_92 ( BL92, BLN92, WL106);
sram_cell_6t_3 inst_cell_106_91 ( BL91, BLN91, WL106);
sram_cell_6t_3 inst_cell_106_90 ( BL90, BLN90, WL106);
sram_cell_6t_3 inst_cell_106_89 ( BL89, BLN89, WL106);
sram_cell_6t_3 inst_cell_106_88 ( BL88, BLN88, WL106);
sram_cell_6t_3 inst_cell_106_87 ( BL87, BLN87, WL106);
sram_cell_6t_3 inst_cell_106_86 ( BL86, BLN86, WL106);
sram_cell_6t_3 inst_cell_106_85 ( BL85, BLN85, WL106);
sram_cell_6t_3 inst_cell_106_84 ( BL84, BLN84, WL106);
sram_cell_6t_3 inst_cell_106_83 ( BL83, BLN83, WL106);
sram_cell_6t_3 inst_cell_106_82 ( BL82, BLN82, WL106);
sram_cell_6t_3 inst_cell_106_81 ( BL81, BLN81, WL106);
sram_cell_6t_3 inst_cell_106_80 ( BL80, BLN80, WL106);
sram_cell_6t_3 inst_cell_106_79 ( BL79, BLN79, WL106);
sram_cell_6t_3 inst_cell_106_78 ( BL78, BLN78, WL106);
sram_cell_6t_3 inst_cell_106_77 ( BL77, BLN77, WL106);
sram_cell_6t_3 inst_cell_106_76 ( BL76, BLN76, WL106);
sram_cell_6t_3 inst_cell_106_75 ( BL75, BLN75, WL106);
sram_cell_6t_3 inst_cell_106_74 ( BL74, BLN74, WL106);
sram_cell_6t_3 inst_cell_106_73 ( BL73, BLN73, WL106);
sram_cell_6t_3 inst_cell_106_72 ( BL72, BLN72, WL106);
sram_cell_6t_3 inst_cell_106_71 ( BL71, BLN71, WL106);
sram_cell_6t_3 inst_cell_106_70 ( BL70, BLN70, WL106);
sram_cell_6t_3 inst_cell_106_69 ( BL69, BLN69, WL106);
sram_cell_6t_3 inst_cell_106_68 ( BL68, BLN68, WL106);
sram_cell_6t_3 inst_cell_106_67 ( BL67, BLN67, WL106);
sram_cell_6t_3 inst_cell_106_66 ( BL66, BLN66, WL106);
sram_cell_6t_3 inst_cell_106_65 ( BL65, BLN65, WL106);
sram_cell_6t_3 inst_cell_106_64 ( BL64, BLN64, WL106);
sram_cell_6t_3 inst_cell_106_63 ( BL63, BLN63, WL106);
sram_cell_6t_3 inst_cell_106_62 ( BL62, BLN62, WL106);
sram_cell_6t_3 inst_cell_106_61 ( BL61, BLN61, WL106);
sram_cell_6t_3 inst_cell_106_60 ( BL60, BLN60, WL106);
sram_cell_6t_3 inst_cell_106_59 ( BL59, BLN59, WL106);
sram_cell_6t_3 inst_cell_106_58 ( BL58, BLN58, WL106);
sram_cell_6t_3 inst_cell_106_57 ( BL57, BLN57, WL106);
sram_cell_6t_3 inst_cell_106_56 ( BL56, BLN56, WL106);
sram_cell_6t_3 inst_cell_106_55 ( BL55, BLN55, WL106);
sram_cell_6t_3 inst_cell_106_54 ( BL54, BLN54, WL106);
sram_cell_6t_3 inst_cell_106_53 ( BL53, BLN53, WL106);
sram_cell_6t_3 inst_cell_106_52 ( BL52, BLN52, WL106);
sram_cell_6t_3 inst_cell_106_51 ( BL51, BLN51, WL106);
sram_cell_6t_3 inst_cell_106_50 ( BL50, BLN50, WL106);
sram_cell_6t_3 inst_cell_106_49 ( BL49, BLN49, WL106);
sram_cell_6t_3 inst_cell_106_48 ( BL48, BLN48, WL106);
sram_cell_6t_3 inst_cell_106_47 ( BL47, BLN47, WL106);
sram_cell_6t_3 inst_cell_106_46 ( BL46, BLN46, WL106);
sram_cell_6t_3 inst_cell_106_45 ( BL45, BLN45, WL106);
sram_cell_6t_3 inst_cell_106_44 ( BL44, BLN44, WL106);
sram_cell_6t_3 inst_cell_106_43 ( BL43, BLN43, WL106);
sram_cell_6t_3 inst_cell_106_42 ( BL42, BLN42, WL106);
sram_cell_6t_3 inst_cell_106_41 ( BL41, BLN41, WL106);
sram_cell_6t_3 inst_cell_106_40 ( BL40, BLN40, WL106);
sram_cell_6t_3 inst_cell_106_39 ( BL39, BLN39, WL106);
sram_cell_6t_3 inst_cell_106_38 ( BL38, BLN38, WL106);
sram_cell_6t_3 inst_cell_106_37 ( BL37, BLN37, WL106);
sram_cell_6t_3 inst_cell_106_36 ( BL36, BLN36, WL106);
sram_cell_6t_3 inst_cell_106_35 ( BL35, BLN35, WL106);
sram_cell_6t_3 inst_cell_106_34 ( BL34, BLN34, WL106);
sram_cell_6t_3 inst_cell_106_33 ( BL33, BLN33, WL106);
sram_cell_6t_3 inst_cell_106_32 ( BL32, BLN32, WL106);
sram_cell_6t_3 inst_cell_106_31 ( BL31, BLN31, WL106);
sram_cell_6t_3 inst_cell_106_30 ( BL30, BLN30, WL106);
sram_cell_6t_3 inst_cell_106_29 ( BL29, BLN29, WL106);
sram_cell_6t_3 inst_cell_106_28 ( BL28, BLN28, WL106);
sram_cell_6t_3 inst_cell_106_27 ( BL27, BLN27, WL106);
sram_cell_6t_3 inst_cell_106_26 ( BL26, BLN26, WL106);
sram_cell_6t_3 inst_cell_106_25 ( BL25, BLN25, WL106);
sram_cell_6t_3 inst_cell_106_24 ( BL24, BLN24, WL106);
sram_cell_6t_3 inst_cell_106_23 ( BL23, BLN23, WL106);
sram_cell_6t_3 inst_cell_106_22 ( BL22, BLN22, WL106);
sram_cell_6t_3 inst_cell_106_21 ( BL21, BLN21, WL106);
sram_cell_6t_3 inst_cell_106_20 ( BL20, BLN20, WL106);
sram_cell_6t_3 inst_cell_106_19 ( BL19, BLN19, WL106);
sram_cell_6t_3 inst_cell_106_18 ( BL18, BLN18, WL106);
sram_cell_6t_3 inst_cell_106_17 ( BL17, BLN17, WL106);
sram_cell_6t_3 inst_cell_106_16 ( BL16, BLN16, WL106);
sram_cell_6t_3 inst_cell_106_15 ( BL15, BLN15, WL106);
sram_cell_6t_3 inst_cell_106_14 ( BL14, BLN14, WL106);
sram_cell_6t_3 inst_cell_106_13 ( BL13, BLN13, WL106);
sram_cell_6t_3 inst_cell_106_12 ( BL12, BLN12, WL106);
sram_cell_6t_3 inst_cell_106_11 ( BL11, BLN11, WL106);
sram_cell_6t_3 inst_cell_106_10 ( BL10, BLN10, WL106);
sram_cell_6t_3 inst_cell_106_9 ( BL9, BLN9, WL106);
sram_cell_6t_3 inst_cell_106_8 ( BL8, BLN8, WL106);
sram_cell_6t_3 inst_cell_106_7 ( BL7, BLN7, WL106);
sram_cell_6t_3 inst_cell_106_6 ( BL6, BLN6, WL106);
sram_cell_6t_3 inst_cell_106_5 ( BL5, BLN5, WL106);
sram_cell_6t_3 inst_cell_106_4 ( BL4, BLN4, WL106);
sram_cell_6t_3 inst_cell_106_3 ( BL3, BLN3, WL106);
sram_cell_6t_3 inst_cell_106_2 ( BL2, BLN2, WL106);
sram_cell_6t_3 inst_cell_106_1 ( BL1, BLN1, WL106);
sram_cell_6t_3 inst_cell_106_0 ( BL0, BLN0, WL106);
sram_cell_6t_3 inst_cell_105_127 ( BL127, BLN127, WL105);
sram_cell_6t_3 inst_cell_105_126 ( BL126, BLN126, WL105);
sram_cell_6t_3 inst_cell_105_125 ( BL125, BLN125, WL105);
sram_cell_6t_3 inst_cell_105_124 ( BL124, BLN124, WL105);
sram_cell_6t_3 inst_cell_105_123 ( BL123, BLN123, WL105);
sram_cell_6t_3 inst_cell_105_122 ( BL122, BLN122, WL105);
sram_cell_6t_3 inst_cell_105_121 ( BL121, BLN121, WL105);
sram_cell_6t_3 inst_cell_105_120 ( BL120, BLN120, WL105);
sram_cell_6t_3 inst_cell_105_119 ( BL119, BLN119, WL105);
sram_cell_6t_3 inst_cell_105_118 ( BL118, BLN118, WL105);
sram_cell_6t_3 inst_cell_105_117 ( BL117, BLN117, WL105);
sram_cell_6t_3 inst_cell_105_116 ( BL116, BLN116, WL105);
sram_cell_6t_3 inst_cell_105_115 ( BL115, BLN115, WL105);
sram_cell_6t_3 inst_cell_105_114 ( BL114, BLN114, WL105);
sram_cell_6t_3 inst_cell_105_113 ( BL113, BLN113, WL105);
sram_cell_6t_3 inst_cell_105_112 ( BL112, BLN112, WL105);
sram_cell_6t_3 inst_cell_105_111 ( BL111, BLN111, WL105);
sram_cell_6t_3 inst_cell_105_110 ( BL110, BLN110, WL105);
sram_cell_6t_3 inst_cell_105_109 ( BL109, BLN109, WL105);
sram_cell_6t_3 inst_cell_105_108 ( BL108, BLN108, WL105);
sram_cell_6t_3 inst_cell_105_107 ( BL107, BLN107, WL105);
sram_cell_6t_3 inst_cell_105_106 ( BL106, BLN106, WL105);
sram_cell_6t_3 inst_cell_105_105 ( BL105, BLN105, WL105);
sram_cell_6t_3 inst_cell_105_104 ( BL104, BLN104, WL105);
sram_cell_6t_3 inst_cell_105_103 ( BL103, BLN103, WL105);
sram_cell_6t_3 inst_cell_105_102 ( BL102, BLN102, WL105);
sram_cell_6t_3 inst_cell_105_101 ( BL101, BLN101, WL105);
sram_cell_6t_3 inst_cell_105_100 ( BL100, BLN100, WL105);
sram_cell_6t_3 inst_cell_105_99 ( BL99, BLN99, WL105);
sram_cell_6t_3 inst_cell_105_98 ( BL98, BLN98, WL105);
sram_cell_6t_3 inst_cell_105_97 ( BL97, BLN97, WL105);
sram_cell_6t_3 inst_cell_105_96 ( BL96, BLN96, WL105);
sram_cell_6t_3 inst_cell_105_95 ( BL95, BLN95, WL105);
sram_cell_6t_3 inst_cell_105_94 ( BL94, BLN94, WL105);
sram_cell_6t_3 inst_cell_105_93 ( BL93, BLN93, WL105);
sram_cell_6t_3 inst_cell_105_92 ( BL92, BLN92, WL105);
sram_cell_6t_3 inst_cell_105_91 ( BL91, BLN91, WL105);
sram_cell_6t_3 inst_cell_105_90 ( BL90, BLN90, WL105);
sram_cell_6t_3 inst_cell_105_89 ( BL89, BLN89, WL105);
sram_cell_6t_3 inst_cell_105_88 ( BL88, BLN88, WL105);
sram_cell_6t_3 inst_cell_105_87 ( BL87, BLN87, WL105);
sram_cell_6t_3 inst_cell_105_86 ( BL86, BLN86, WL105);
sram_cell_6t_3 inst_cell_105_85 ( BL85, BLN85, WL105);
sram_cell_6t_3 inst_cell_105_84 ( BL84, BLN84, WL105);
sram_cell_6t_3 inst_cell_105_83 ( BL83, BLN83, WL105);
sram_cell_6t_3 inst_cell_105_82 ( BL82, BLN82, WL105);
sram_cell_6t_3 inst_cell_105_81 ( BL81, BLN81, WL105);
sram_cell_6t_3 inst_cell_105_80 ( BL80, BLN80, WL105);
sram_cell_6t_3 inst_cell_105_79 ( BL79, BLN79, WL105);
sram_cell_6t_3 inst_cell_105_78 ( BL78, BLN78, WL105);
sram_cell_6t_3 inst_cell_105_77 ( BL77, BLN77, WL105);
sram_cell_6t_3 inst_cell_105_76 ( BL76, BLN76, WL105);
sram_cell_6t_3 inst_cell_105_75 ( BL75, BLN75, WL105);
sram_cell_6t_3 inst_cell_105_74 ( BL74, BLN74, WL105);
sram_cell_6t_3 inst_cell_105_73 ( BL73, BLN73, WL105);
sram_cell_6t_3 inst_cell_105_72 ( BL72, BLN72, WL105);
sram_cell_6t_3 inst_cell_105_71 ( BL71, BLN71, WL105);
sram_cell_6t_3 inst_cell_105_70 ( BL70, BLN70, WL105);
sram_cell_6t_3 inst_cell_105_69 ( BL69, BLN69, WL105);
sram_cell_6t_3 inst_cell_105_68 ( BL68, BLN68, WL105);
sram_cell_6t_3 inst_cell_105_67 ( BL67, BLN67, WL105);
sram_cell_6t_3 inst_cell_105_66 ( BL66, BLN66, WL105);
sram_cell_6t_3 inst_cell_105_65 ( BL65, BLN65, WL105);
sram_cell_6t_3 inst_cell_105_64 ( BL64, BLN64, WL105);
sram_cell_6t_3 inst_cell_105_63 ( BL63, BLN63, WL105);
sram_cell_6t_3 inst_cell_105_62 ( BL62, BLN62, WL105);
sram_cell_6t_3 inst_cell_105_61 ( BL61, BLN61, WL105);
sram_cell_6t_3 inst_cell_105_60 ( BL60, BLN60, WL105);
sram_cell_6t_3 inst_cell_105_59 ( BL59, BLN59, WL105);
sram_cell_6t_3 inst_cell_105_58 ( BL58, BLN58, WL105);
sram_cell_6t_3 inst_cell_105_57 ( BL57, BLN57, WL105);
sram_cell_6t_3 inst_cell_105_56 ( BL56, BLN56, WL105);
sram_cell_6t_3 inst_cell_105_55 ( BL55, BLN55, WL105);
sram_cell_6t_3 inst_cell_105_54 ( BL54, BLN54, WL105);
sram_cell_6t_3 inst_cell_105_53 ( BL53, BLN53, WL105);
sram_cell_6t_3 inst_cell_105_52 ( BL52, BLN52, WL105);
sram_cell_6t_3 inst_cell_105_51 ( BL51, BLN51, WL105);
sram_cell_6t_3 inst_cell_105_50 ( BL50, BLN50, WL105);
sram_cell_6t_3 inst_cell_105_49 ( BL49, BLN49, WL105);
sram_cell_6t_3 inst_cell_105_48 ( BL48, BLN48, WL105);
sram_cell_6t_3 inst_cell_105_47 ( BL47, BLN47, WL105);
sram_cell_6t_3 inst_cell_105_46 ( BL46, BLN46, WL105);
sram_cell_6t_3 inst_cell_105_45 ( BL45, BLN45, WL105);
sram_cell_6t_3 inst_cell_105_44 ( BL44, BLN44, WL105);
sram_cell_6t_3 inst_cell_105_43 ( BL43, BLN43, WL105);
sram_cell_6t_3 inst_cell_105_42 ( BL42, BLN42, WL105);
sram_cell_6t_3 inst_cell_105_41 ( BL41, BLN41, WL105);
sram_cell_6t_3 inst_cell_105_40 ( BL40, BLN40, WL105);
sram_cell_6t_3 inst_cell_105_39 ( BL39, BLN39, WL105);
sram_cell_6t_3 inst_cell_105_38 ( BL38, BLN38, WL105);
sram_cell_6t_3 inst_cell_105_37 ( BL37, BLN37, WL105);
sram_cell_6t_3 inst_cell_105_36 ( BL36, BLN36, WL105);
sram_cell_6t_3 inst_cell_105_35 ( BL35, BLN35, WL105);
sram_cell_6t_3 inst_cell_105_34 ( BL34, BLN34, WL105);
sram_cell_6t_3 inst_cell_105_33 ( BL33, BLN33, WL105);
sram_cell_6t_3 inst_cell_105_32 ( BL32, BLN32, WL105);
sram_cell_6t_3 inst_cell_105_31 ( BL31, BLN31, WL105);
sram_cell_6t_3 inst_cell_105_30 ( BL30, BLN30, WL105);
sram_cell_6t_3 inst_cell_105_29 ( BL29, BLN29, WL105);
sram_cell_6t_3 inst_cell_105_28 ( BL28, BLN28, WL105);
sram_cell_6t_3 inst_cell_105_27 ( BL27, BLN27, WL105);
sram_cell_6t_3 inst_cell_105_26 ( BL26, BLN26, WL105);
sram_cell_6t_3 inst_cell_105_25 ( BL25, BLN25, WL105);
sram_cell_6t_3 inst_cell_105_24 ( BL24, BLN24, WL105);
sram_cell_6t_3 inst_cell_105_23 ( BL23, BLN23, WL105);
sram_cell_6t_3 inst_cell_105_22 ( BL22, BLN22, WL105);
sram_cell_6t_3 inst_cell_105_21 ( BL21, BLN21, WL105);
sram_cell_6t_3 inst_cell_105_20 ( BL20, BLN20, WL105);
sram_cell_6t_3 inst_cell_105_19 ( BL19, BLN19, WL105);
sram_cell_6t_3 inst_cell_105_18 ( BL18, BLN18, WL105);
sram_cell_6t_3 inst_cell_105_17 ( BL17, BLN17, WL105);
sram_cell_6t_3 inst_cell_105_16 ( BL16, BLN16, WL105);
sram_cell_6t_3 inst_cell_105_15 ( BL15, BLN15, WL105);
sram_cell_6t_3 inst_cell_105_14 ( BL14, BLN14, WL105);
sram_cell_6t_3 inst_cell_105_13 ( BL13, BLN13, WL105);
sram_cell_6t_3 inst_cell_105_12 ( BL12, BLN12, WL105);
sram_cell_6t_3 inst_cell_105_11 ( BL11, BLN11, WL105);
sram_cell_6t_3 inst_cell_105_10 ( BL10, BLN10, WL105);
sram_cell_6t_3 inst_cell_105_9 ( BL9, BLN9, WL105);
sram_cell_6t_3 inst_cell_105_8 ( BL8, BLN8, WL105);
sram_cell_6t_3 inst_cell_105_7 ( BL7, BLN7, WL105);
sram_cell_6t_3 inst_cell_105_6 ( BL6, BLN6, WL105);
sram_cell_6t_3 inst_cell_105_5 ( BL5, BLN5, WL105);
sram_cell_6t_3 inst_cell_105_4 ( BL4, BLN4, WL105);
sram_cell_6t_3 inst_cell_105_3 ( BL3, BLN3, WL105);
sram_cell_6t_3 inst_cell_105_2 ( BL2, BLN2, WL105);
sram_cell_6t_3 inst_cell_105_1 ( BL1, BLN1, WL105);
sram_cell_6t_3 inst_cell_105_0 ( BL0, BLN0, WL105);
sram_cell_6t_3 inst_cell_104_127 ( BL127, BLN127, WL104);
sram_cell_6t_3 inst_cell_104_126 ( BL126, BLN126, WL104);
sram_cell_6t_3 inst_cell_104_125 ( BL125, BLN125, WL104);
sram_cell_6t_3 inst_cell_104_124 ( BL124, BLN124, WL104);
sram_cell_6t_3 inst_cell_104_123 ( BL123, BLN123, WL104);
sram_cell_6t_3 inst_cell_104_122 ( BL122, BLN122, WL104);
sram_cell_6t_3 inst_cell_104_121 ( BL121, BLN121, WL104);
sram_cell_6t_3 inst_cell_104_120 ( BL120, BLN120, WL104);
sram_cell_6t_3 inst_cell_104_119 ( BL119, BLN119, WL104);
sram_cell_6t_3 inst_cell_104_118 ( BL118, BLN118, WL104);
sram_cell_6t_3 inst_cell_104_117 ( BL117, BLN117, WL104);
sram_cell_6t_3 inst_cell_104_116 ( BL116, BLN116, WL104);
sram_cell_6t_3 inst_cell_104_115 ( BL115, BLN115, WL104);
sram_cell_6t_3 inst_cell_104_114 ( BL114, BLN114, WL104);
sram_cell_6t_3 inst_cell_104_113 ( BL113, BLN113, WL104);
sram_cell_6t_3 inst_cell_104_112 ( BL112, BLN112, WL104);
sram_cell_6t_3 inst_cell_104_111 ( BL111, BLN111, WL104);
sram_cell_6t_3 inst_cell_104_110 ( BL110, BLN110, WL104);
sram_cell_6t_3 inst_cell_104_109 ( BL109, BLN109, WL104);
sram_cell_6t_3 inst_cell_104_108 ( BL108, BLN108, WL104);
sram_cell_6t_3 inst_cell_104_107 ( BL107, BLN107, WL104);
sram_cell_6t_3 inst_cell_104_106 ( BL106, BLN106, WL104);
sram_cell_6t_3 inst_cell_104_105 ( BL105, BLN105, WL104);
sram_cell_6t_3 inst_cell_104_104 ( BL104, BLN104, WL104);
sram_cell_6t_3 inst_cell_104_103 ( BL103, BLN103, WL104);
sram_cell_6t_3 inst_cell_104_102 ( BL102, BLN102, WL104);
sram_cell_6t_3 inst_cell_104_101 ( BL101, BLN101, WL104);
sram_cell_6t_3 inst_cell_104_100 ( BL100, BLN100, WL104);
sram_cell_6t_3 inst_cell_104_99 ( BL99, BLN99, WL104);
sram_cell_6t_3 inst_cell_104_98 ( BL98, BLN98, WL104);
sram_cell_6t_3 inst_cell_104_97 ( BL97, BLN97, WL104);
sram_cell_6t_3 inst_cell_104_96 ( BL96, BLN96, WL104);
sram_cell_6t_3 inst_cell_104_95 ( BL95, BLN95, WL104);
sram_cell_6t_3 inst_cell_104_94 ( BL94, BLN94, WL104);
sram_cell_6t_3 inst_cell_104_93 ( BL93, BLN93, WL104);
sram_cell_6t_3 inst_cell_104_92 ( BL92, BLN92, WL104);
sram_cell_6t_3 inst_cell_104_91 ( BL91, BLN91, WL104);
sram_cell_6t_3 inst_cell_104_90 ( BL90, BLN90, WL104);
sram_cell_6t_3 inst_cell_104_89 ( BL89, BLN89, WL104);
sram_cell_6t_3 inst_cell_104_88 ( BL88, BLN88, WL104);
sram_cell_6t_3 inst_cell_104_87 ( BL87, BLN87, WL104);
sram_cell_6t_3 inst_cell_104_86 ( BL86, BLN86, WL104);
sram_cell_6t_3 inst_cell_104_85 ( BL85, BLN85, WL104);
sram_cell_6t_3 inst_cell_104_84 ( BL84, BLN84, WL104);
sram_cell_6t_3 inst_cell_104_83 ( BL83, BLN83, WL104);
sram_cell_6t_3 inst_cell_104_82 ( BL82, BLN82, WL104);
sram_cell_6t_3 inst_cell_104_81 ( BL81, BLN81, WL104);
sram_cell_6t_3 inst_cell_104_80 ( BL80, BLN80, WL104);
sram_cell_6t_3 inst_cell_104_79 ( BL79, BLN79, WL104);
sram_cell_6t_3 inst_cell_104_78 ( BL78, BLN78, WL104);
sram_cell_6t_3 inst_cell_104_77 ( BL77, BLN77, WL104);
sram_cell_6t_3 inst_cell_104_76 ( BL76, BLN76, WL104);
sram_cell_6t_3 inst_cell_104_75 ( BL75, BLN75, WL104);
sram_cell_6t_3 inst_cell_104_74 ( BL74, BLN74, WL104);
sram_cell_6t_3 inst_cell_104_73 ( BL73, BLN73, WL104);
sram_cell_6t_3 inst_cell_104_72 ( BL72, BLN72, WL104);
sram_cell_6t_3 inst_cell_104_71 ( BL71, BLN71, WL104);
sram_cell_6t_3 inst_cell_104_70 ( BL70, BLN70, WL104);
sram_cell_6t_3 inst_cell_104_69 ( BL69, BLN69, WL104);
sram_cell_6t_3 inst_cell_104_68 ( BL68, BLN68, WL104);
sram_cell_6t_3 inst_cell_104_67 ( BL67, BLN67, WL104);
sram_cell_6t_3 inst_cell_104_66 ( BL66, BLN66, WL104);
sram_cell_6t_3 inst_cell_104_65 ( BL65, BLN65, WL104);
sram_cell_6t_3 inst_cell_104_64 ( BL64, BLN64, WL104);
sram_cell_6t_3 inst_cell_104_63 ( BL63, BLN63, WL104);
sram_cell_6t_3 inst_cell_104_62 ( BL62, BLN62, WL104);
sram_cell_6t_3 inst_cell_104_61 ( BL61, BLN61, WL104);
sram_cell_6t_3 inst_cell_104_60 ( BL60, BLN60, WL104);
sram_cell_6t_3 inst_cell_104_59 ( BL59, BLN59, WL104);
sram_cell_6t_3 inst_cell_104_58 ( BL58, BLN58, WL104);
sram_cell_6t_3 inst_cell_104_57 ( BL57, BLN57, WL104);
sram_cell_6t_3 inst_cell_104_56 ( BL56, BLN56, WL104);
sram_cell_6t_3 inst_cell_104_55 ( BL55, BLN55, WL104);
sram_cell_6t_3 inst_cell_104_54 ( BL54, BLN54, WL104);
sram_cell_6t_3 inst_cell_104_53 ( BL53, BLN53, WL104);
sram_cell_6t_3 inst_cell_104_52 ( BL52, BLN52, WL104);
sram_cell_6t_3 inst_cell_104_51 ( BL51, BLN51, WL104);
sram_cell_6t_3 inst_cell_104_50 ( BL50, BLN50, WL104);
sram_cell_6t_3 inst_cell_104_49 ( BL49, BLN49, WL104);
sram_cell_6t_3 inst_cell_104_48 ( BL48, BLN48, WL104);
sram_cell_6t_3 inst_cell_104_47 ( BL47, BLN47, WL104);
sram_cell_6t_3 inst_cell_104_46 ( BL46, BLN46, WL104);
sram_cell_6t_3 inst_cell_104_45 ( BL45, BLN45, WL104);
sram_cell_6t_3 inst_cell_104_44 ( BL44, BLN44, WL104);
sram_cell_6t_3 inst_cell_104_43 ( BL43, BLN43, WL104);
sram_cell_6t_3 inst_cell_104_42 ( BL42, BLN42, WL104);
sram_cell_6t_3 inst_cell_104_41 ( BL41, BLN41, WL104);
sram_cell_6t_3 inst_cell_104_40 ( BL40, BLN40, WL104);
sram_cell_6t_3 inst_cell_104_39 ( BL39, BLN39, WL104);
sram_cell_6t_3 inst_cell_104_38 ( BL38, BLN38, WL104);
sram_cell_6t_3 inst_cell_104_37 ( BL37, BLN37, WL104);
sram_cell_6t_3 inst_cell_104_36 ( BL36, BLN36, WL104);
sram_cell_6t_3 inst_cell_104_35 ( BL35, BLN35, WL104);
sram_cell_6t_3 inst_cell_104_34 ( BL34, BLN34, WL104);
sram_cell_6t_3 inst_cell_104_33 ( BL33, BLN33, WL104);
sram_cell_6t_3 inst_cell_104_32 ( BL32, BLN32, WL104);
sram_cell_6t_3 inst_cell_104_31 ( BL31, BLN31, WL104);
sram_cell_6t_3 inst_cell_104_30 ( BL30, BLN30, WL104);
sram_cell_6t_3 inst_cell_104_29 ( BL29, BLN29, WL104);
sram_cell_6t_3 inst_cell_104_28 ( BL28, BLN28, WL104);
sram_cell_6t_3 inst_cell_104_27 ( BL27, BLN27, WL104);
sram_cell_6t_3 inst_cell_104_26 ( BL26, BLN26, WL104);
sram_cell_6t_3 inst_cell_104_25 ( BL25, BLN25, WL104);
sram_cell_6t_3 inst_cell_104_24 ( BL24, BLN24, WL104);
sram_cell_6t_3 inst_cell_104_23 ( BL23, BLN23, WL104);
sram_cell_6t_3 inst_cell_104_22 ( BL22, BLN22, WL104);
sram_cell_6t_3 inst_cell_104_21 ( BL21, BLN21, WL104);
sram_cell_6t_3 inst_cell_104_20 ( BL20, BLN20, WL104);
sram_cell_6t_3 inst_cell_104_19 ( BL19, BLN19, WL104);
sram_cell_6t_3 inst_cell_104_18 ( BL18, BLN18, WL104);
sram_cell_6t_3 inst_cell_104_17 ( BL17, BLN17, WL104);
sram_cell_6t_3 inst_cell_104_16 ( BL16, BLN16, WL104);
sram_cell_6t_3 inst_cell_104_15 ( BL15, BLN15, WL104);
sram_cell_6t_3 inst_cell_104_14 ( BL14, BLN14, WL104);
sram_cell_6t_3 inst_cell_104_13 ( BL13, BLN13, WL104);
sram_cell_6t_3 inst_cell_104_12 ( BL12, BLN12, WL104);
sram_cell_6t_3 inst_cell_104_11 ( BL11, BLN11, WL104);
sram_cell_6t_3 inst_cell_104_10 ( BL10, BLN10, WL104);
sram_cell_6t_3 inst_cell_104_9 ( BL9, BLN9, WL104);
sram_cell_6t_3 inst_cell_104_8 ( BL8, BLN8, WL104);
sram_cell_6t_3 inst_cell_104_7 ( BL7, BLN7, WL104);
sram_cell_6t_3 inst_cell_104_6 ( BL6, BLN6, WL104);
sram_cell_6t_3 inst_cell_104_5 ( BL5, BLN5, WL104);
sram_cell_6t_3 inst_cell_104_4 ( BL4, BLN4, WL104);
sram_cell_6t_3 inst_cell_104_3 ( BL3, BLN3, WL104);
sram_cell_6t_3 inst_cell_104_2 ( BL2, BLN2, WL104);
sram_cell_6t_3 inst_cell_104_1 ( BL1, BLN1, WL104);
sram_cell_6t_3 inst_cell_104_0 ( BL0, BLN0, WL104);
sram_cell_6t_3 inst_cell_103_127 ( BL127, BLN127, WL103);
sram_cell_6t_3 inst_cell_103_126 ( BL126, BLN126, WL103);
sram_cell_6t_3 inst_cell_103_125 ( BL125, BLN125, WL103);
sram_cell_6t_3 inst_cell_103_124 ( BL124, BLN124, WL103);
sram_cell_6t_3 inst_cell_103_123 ( BL123, BLN123, WL103);
sram_cell_6t_3 inst_cell_103_122 ( BL122, BLN122, WL103);
sram_cell_6t_3 inst_cell_103_121 ( BL121, BLN121, WL103);
sram_cell_6t_3 inst_cell_103_120 ( BL120, BLN120, WL103);
sram_cell_6t_3 inst_cell_103_119 ( BL119, BLN119, WL103);
sram_cell_6t_3 inst_cell_103_118 ( BL118, BLN118, WL103);
sram_cell_6t_3 inst_cell_103_117 ( BL117, BLN117, WL103);
sram_cell_6t_3 inst_cell_103_116 ( BL116, BLN116, WL103);
sram_cell_6t_3 inst_cell_103_115 ( BL115, BLN115, WL103);
sram_cell_6t_3 inst_cell_103_114 ( BL114, BLN114, WL103);
sram_cell_6t_3 inst_cell_103_113 ( BL113, BLN113, WL103);
sram_cell_6t_3 inst_cell_103_112 ( BL112, BLN112, WL103);
sram_cell_6t_3 inst_cell_103_111 ( BL111, BLN111, WL103);
sram_cell_6t_3 inst_cell_103_110 ( BL110, BLN110, WL103);
sram_cell_6t_3 inst_cell_103_109 ( BL109, BLN109, WL103);
sram_cell_6t_3 inst_cell_103_108 ( BL108, BLN108, WL103);
sram_cell_6t_3 inst_cell_103_107 ( BL107, BLN107, WL103);
sram_cell_6t_3 inst_cell_103_106 ( BL106, BLN106, WL103);
sram_cell_6t_3 inst_cell_103_105 ( BL105, BLN105, WL103);
sram_cell_6t_3 inst_cell_103_104 ( BL104, BLN104, WL103);
sram_cell_6t_3 inst_cell_103_103 ( BL103, BLN103, WL103);
sram_cell_6t_3 inst_cell_103_102 ( BL102, BLN102, WL103);
sram_cell_6t_3 inst_cell_103_101 ( BL101, BLN101, WL103);
sram_cell_6t_3 inst_cell_103_100 ( BL100, BLN100, WL103);
sram_cell_6t_3 inst_cell_103_99 ( BL99, BLN99, WL103);
sram_cell_6t_3 inst_cell_103_98 ( BL98, BLN98, WL103);
sram_cell_6t_3 inst_cell_103_97 ( BL97, BLN97, WL103);
sram_cell_6t_3 inst_cell_103_96 ( BL96, BLN96, WL103);
sram_cell_6t_3 inst_cell_103_95 ( BL95, BLN95, WL103);
sram_cell_6t_3 inst_cell_103_94 ( BL94, BLN94, WL103);
sram_cell_6t_3 inst_cell_103_93 ( BL93, BLN93, WL103);
sram_cell_6t_3 inst_cell_103_92 ( BL92, BLN92, WL103);
sram_cell_6t_3 inst_cell_103_91 ( BL91, BLN91, WL103);
sram_cell_6t_3 inst_cell_103_90 ( BL90, BLN90, WL103);
sram_cell_6t_3 inst_cell_103_89 ( BL89, BLN89, WL103);
sram_cell_6t_3 inst_cell_103_88 ( BL88, BLN88, WL103);
sram_cell_6t_3 inst_cell_103_87 ( BL87, BLN87, WL103);
sram_cell_6t_3 inst_cell_103_86 ( BL86, BLN86, WL103);
sram_cell_6t_3 inst_cell_103_85 ( BL85, BLN85, WL103);
sram_cell_6t_3 inst_cell_103_84 ( BL84, BLN84, WL103);
sram_cell_6t_3 inst_cell_103_83 ( BL83, BLN83, WL103);
sram_cell_6t_3 inst_cell_103_82 ( BL82, BLN82, WL103);
sram_cell_6t_3 inst_cell_103_81 ( BL81, BLN81, WL103);
sram_cell_6t_3 inst_cell_103_80 ( BL80, BLN80, WL103);
sram_cell_6t_3 inst_cell_103_79 ( BL79, BLN79, WL103);
sram_cell_6t_3 inst_cell_103_78 ( BL78, BLN78, WL103);
sram_cell_6t_3 inst_cell_103_77 ( BL77, BLN77, WL103);
sram_cell_6t_3 inst_cell_103_76 ( BL76, BLN76, WL103);
sram_cell_6t_3 inst_cell_103_75 ( BL75, BLN75, WL103);
sram_cell_6t_3 inst_cell_103_74 ( BL74, BLN74, WL103);
sram_cell_6t_3 inst_cell_103_73 ( BL73, BLN73, WL103);
sram_cell_6t_3 inst_cell_103_72 ( BL72, BLN72, WL103);
sram_cell_6t_3 inst_cell_103_71 ( BL71, BLN71, WL103);
sram_cell_6t_3 inst_cell_103_70 ( BL70, BLN70, WL103);
sram_cell_6t_3 inst_cell_103_69 ( BL69, BLN69, WL103);
sram_cell_6t_3 inst_cell_103_68 ( BL68, BLN68, WL103);
sram_cell_6t_3 inst_cell_103_67 ( BL67, BLN67, WL103);
sram_cell_6t_3 inst_cell_103_66 ( BL66, BLN66, WL103);
sram_cell_6t_3 inst_cell_103_65 ( BL65, BLN65, WL103);
sram_cell_6t_3 inst_cell_103_64 ( BL64, BLN64, WL103);
sram_cell_6t_3 inst_cell_103_63 ( BL63, BLN63, WL103);
sram_cell_6t_3 inst_cell_103_62 ( BL62, BLN62, WL103);
sram_cell_6t_3 inst_cell_103_61 ( BL61, BLN61, WL103);
sram_cell_6t_3 inst_cell_103_60 ( BL60, BLN60, WL103);
sram_cell_6t_3 inst_cell_103_59 ( BL59, BLN59, WL103);
sram_cell_6t_3 inst_cell_103_58 ( BL58, BLN58, WL103);
sram_cell_6t_3 inst_cell_103_57 ( BL57, BLN57, WL103);
sram_cell_6t_3 inst_cell_103_56 ( BL56, BLN56, WL103);
sram_cell_6t_3 inst_cell_103_55 ( BL55, BLN55, WL103);
sram_cell_6t_3 inst_cell_103_54 ( BL54, BLN54, WL103);
sram_cell_6t_3 inst_cell_103_53 ( BL53, BLN53, WL103);
sram_cell_6t_3 inst_cell_103_52 ( BL52, BLN52, WL103);
sram_cell_6t_3 inst_cell_103_51 ( BL51, BLN51, WL103);
sram_cell_6t_3 inst_cell_103_50 ( BL50, BLN50, WL103);
sram_cell_6t_3 inst_cell_103_49 ( BL49, BLN49, WL103);
sram_cell_6t_3 inst_cell_103_48 ( BL48, BLN48, WL103);
sram_cell_6t_3 inst_cell_103_47 ( BL47, BLN47, WL103);
sram_cell_6t_3 inst_cell_103_46 ( BL46, BLN46, WL103);
sram_cell_6t_3 inst_cell_103_45 ( BL45, BLN45, WL103);
sram_cell_6t_3 inst_cell_103_44 ( BL44, BLN44, WL103);
sram_cell_6t_3 inst_cell_103_43 ( BL43, BLN43, WL103);
sram_cell_6t_3 inst_cell_103_42 ( BL42, BLN42, WL103);
sram_cell_6t_3 inst_cell_103_41 ( BL41, BLN41, WL103);
sram_cell_6t_3 inst_cell_103_40 ( BL40, BLN40, WL103);
sram_cell_6t_3 inst_cell_103_39 ( BL39, BLN39, WL103);
sram_cell_6t_3 inst_cell_103_38 ( BL38, BLN38, WL103);
sram_cell_6t_3 inst_cell_103_37 ( BL37, BLN37, WL103);
sram_cell_6t_3 inst_cell_103_36 ( BL36, BLN36, WL103);
sram_cell_6t_3 inst_cell_103_35 ( BL35, BLN35, WL103);
sram_cell_6t_3 inst_cell_103_34 ( BL34, BLN34, WL103);
sram_cell_6t_3 inst_cell_103_33 ( BL33, BLN33, WL103);
sram_cell_6t_3 inst_cell_103_32 ( BL32, BLN32, WL103);
sram_cell_6t_3 inst_cell_103_31 ( BL31, BLN31, WL103);
sram_cell_6t_3 inst_cell_103_30 ( BL30, BLN30, WL103);
sram_cell_6t_3 inst_cell_103_29 ( BL29, BLN29, WL103);
sram_cell_6t_3 inst_cell_103_28 ( BL28, BLN28, WL103);
sram_cell_6t_3 inst_cell_103_27 ( BL27, BLN27, WL103);
sram_cell_6t_3 inst_cell_103_26 ( BL26, BLN26, WL103);
sram_cell_6t_3 inst_cell_103_25 ( BL25, BLN25, WL103);
sram_cell_6t_3 inst_cell_103_24 ( BL24, BLN24, WL103);
sram_cell_6t_3 inst_cell_103_23 ( BL23, BLN23, WL103);
sram_cell_6t_3 inst_cell_103_22 ( BL22, BLN22, WL103);
sram_cell_6t_3 inst_cell_103_21 ( BL21, BLN21, WL103);
sram_cell_6t_3 inst_cell_103_20 ( BL20, BLN20, WL103);
sram_cell_6t_3 inst_cell_103_19 ( BL19, BLN19, WL103);
sram_cell_6t_3 inst_cell_103_18 ( BL18, BLN18, WL103);
sram_cell_6t_3 inst_cell_103_17 ( BL17, BLN17, WL103);
sram_cell_6t_3 inst_cell_103_16 ( BL16, BLN16, WL103);
sram_cell_6t_3 inst_cell_103_15 ( BL15, BLN15, WL103);
sram_cell_6t_3 inst_cell_103_14 ( BL14, BLN14, WL103);
sram_cell_6t_3 inst_cell_103_13 ( BL13, BLN13, WL103);
sram_cell_6t_3 inst_cell_103_12 ( BL12, BLN12, WL103);
sram_cell_6t_3 inst_cell_103_11 ( BL11, BLN11, WL103);
sram_cell_6t_3 inst_cell_103_10 ( BL10, BLN10, WL103);
sram_cell_6t_3 inst_cell_103_9 ( BL9, BLN9, WL103);
sram_cell_6t_3 inst_cell_103_8 ( BL8, BLN8, WL103);
sram_cell_6t_3 inst_cell_103_7 ( BL7, BLN7, WL103);
sram_cell_6t_3 inst_cell_103_6 ( BL6, BLN6, WL103);
sram_cell_6t_3 inst_cell_103_5 ( BL5, BLN5, WL103);
sram_cell_6t_3 inst_cell_103_4 ( BL4, BLN4, WL103);
sram_cell_6t_3 inst_cell_103_3 ( BL3, BLN3, WL103);
sram_cell_6t_3 inst_cell_103_2 ( BL2, BLN2, WL103);
sram_cell_6t_3 inst_cell_103_1 ( BL1, BLN1, WL103);
sram_cell_6t_3 inst_cell_103_0 ( BL0, BLN0, WL103);
sram_cell_6t_3 inst_cell_102_127 ( BL127, BLN127, WL102);
sram_cell_6t_3 inst_cell_102_126 ( BL126, BLN126, WL102);
sram_cell_6t_3 inst_cell_102_125 ( BL125, BLN125, WL102);
sram_cell_6t_3 inst_cell_102_124 ( BL124, BLN124, WL102);
sram_cell_6t_3 inst_cell_102_123 ( BL123, BLN123, WL102);
sram_cell_6t_3 inst_cell_102_122 ( BL122, BLN122, WL102);
sram_cell_6t_3 inst_cell_102_121 ( BL121, BLN121, WL102);
sram_cell_6t_3 inst_cell_102_120 ( BL120, BLN120, WL102);
sram_cell_6t_3 inst_cell_102_119 ( BL119, BLN119, WL102);
sram_cell_6t_3 inst_cell_102_118 ( BL118, BLN118, WL102);
sram_cell_6t_3 inst_cell_102_117 ( BL117, BLN117, WL102);
sram_cell_6t_3 inst_cell_102_116 ( BL116, BLN116, WL102);
sram_cell_6t_3 inst_cell_102_115 ( BL115, BLN115, WL102);
sram_cell_6t_3 inst_cell_102_114 ( BL114, BLN114, WL102);
sram_cell_6t_3 inst_cell_102_113 ( BL113, BLN113, WL102);
sram_cell_6t_3 inst_cell_102_112 ( BL112, BLN112, WL102);
sram_cell_6t_3 inst_cell_102_111 ( BL111, BLN111, WL102);
sram_cell_6t_3 inst_cell_102_110 ( BL110, BLN110, WL102);
sram_cell_6t_3 inst_cell_102_109 ( BL109, BLN109, WL102);
sram_cell_6t_3 inst_cell_102_108 ( BL108, BLN108, WL102);
sram_cell_6t_3 inst_cell_102_107 ( BL107, BLN107, WL102);
sram_cell_6t_3 inst_cell_102_106 ( BL106, BLN106, WL102);
sram_cell_6t_3 inst_cell_102_105 ( BL105, BLN105, WL102);
sram_cell_6t_3 inst_cell_102_104 ( BL104, BLN104, WL102);
sram_cell_6t_3 inst_cell_102_103 ( BL103, BLN103, WL102);
sram_cell_6t_3 inst_cell_102_102 ( BL102, BLN102, WL102);
sram_cell_6t_3 inst_cell_102_101 ( BL101, BLN101, WL102);
sram_cell_6t_3 inst_cell_102_100 ( BL100, BLN100, WL102);
sram_cell_6t_3 inst_cell_102_99 ( BL99, BLN99, WL102);
sram_cell_6t_3 inst_cell_102_98 ( BL98, BLN98, WL102);
sram_cell_6t_3 inst_cell_102_97 ( BL97, BLN97, WL102);
sram_cell_6t_3 inst_cell_102_96 ( BL96, BLN96, WL102);
sram_cell_6t_3 inst_cell_102_95 ( BL95, BLN95, WL102);
sram_cell_6t_3 inst_cell_102_94 ( BL94, BLN94, WL102);
sram_cell_6t_3 inst_cell_102_93 ( BL93, BLN93, WL102);
sram_cell_6t_3 inst_cell_102_92 ( BL92, BLN92, WL102);
sram_cell_6t_3 inst_cell_102_91 ( BL91, BLN91, WL102);
sram_cell_6t_3 inst_cell_102_90 ( BL90, BLN90, WL102);
sram_cell_6t_3 inst_cell_102_89 ( BL89, BLN89, WL102);
sram_cell_6t_3 inst_cell_102_88 ( BL88, BLN88, WL102);
sram_cell_6t_3 inst_cell_102_87 ( BL87, BLN87, WL102);
sram_cell_6t_3 inst_cell_102_86 ( BL86, BLN86, WL102);
sram_cell_6t_3 inst_cell_102_85 ( BL85, BLN85, WL102);
sram_cell_6t_3 inst_cell_102_84 ( BL84, BLN84, WL102);
sram_cell_6t_3 inst_cell_102_83 ( BL83, BLN83, WL102);
sram_cell_6t_3 inst_cell_102_82 ( BL82, BLN82, WL102);
sram_cell_6t_3 inst_cell_102_81 ( BL81, BLN81, WL102);
sram_cell_6t_3 inst_cell_102_80 ( BL80, BLN80, WL102);
sram_cell_6t_3 inst_cell_102_79 ( BL79, BLN79, WL102);
sram_cell_6t_3 inst_cell_102_78 ( BL78, BLN78, WL102);
sram_cell_6t_3 inst_cell_102_77 ( BL77, BLN77, WL102);
sram_cell_6t_3 inst_cell_102_76 ( BL76, BLN76, WL102);
sram_cell_6t_3 inst_cell_102_75 ( BL75, BLN75, WL102);
sram_cell_6t_3 inst_cell_102_74 ( BL74, BLN74, WL102);
sram_cell_6t_3 inst_cell_102_73 ( BL73, BLN73, WL102);
sram_cell_6t_3 inst_cell_102_72 ( BL72, BLN72, WL102);
sram_cell_6t_3 inst_cell_102_71 ( BL71, BLN71, WL102);
sram_cell_6t_3 inst_cell_102_70 ( BL70, BLN70, WL102);
sram_cell_6t_3 inst_cell_102_69 ( BL69, BLN69, WL102);
sram_cell_6t_3 inst_cell_102_68 ( BL68, BLN68, WL102);
sram_cell_6t_3 inst_cell_102_67 ( BL67, BLN67, WL102);
sram_cell_6t_3 inst_cell_102_66 ( BL66, BLN66, WL102);
sram_cell_6t_3 inst_cell_102_65 ( BL65, BLN65, WL102);
sram_cell_6t_3 inst_cell_102_64 ( BL64, BLN64, WL102);
sram_cell_6t_3 inst_cell_102_63 ( BL63, BLN63, WL102);
sram_cell_6t_3 inst_cell_102_62 ( BL62, BLN62, WL102);
sram_cell_6t_3 inst_cell_102_61 ( BL61, BLN61, WL102);
sram_cell_6t_3 inst_cell_102_60 ( BL60, BLN60, WL102);
sram_cell_6t_3 inst_cell_102_59 ( BL59, BLN59, WL102);
sram_cell_6t_3 inst_cell_102_58 ( BL58, BLN58, WL102);
sram_cell_6t_3 inst_cell_102_57 ( BL57, BLN57, WL102);
sram_cell_6t_3 inst_cell_102_56 ( BL56, BLN56, WL102);
sram_cell_6t_3 inst_cell_102_55 ( BL55, BLN55, WL102);
sram_cell_6t_3 inst_cell_102_54 ( BL54, BLN54, WL102);
sram_cell_6t_3 inst_cell_102_53 ( BL53, BLN53, WL102);
sram_cell_6t_3 inst_cell_102_52 ( BL52, BLN52, WL102);
sram_cell_6t_3 inst_cell_102_51 ( BL51, BLN51, WL102);
sram_cell_6t_3 inst_cell_102_50 ( BL50, BLN50, WL102);
sram_cell_6t_3 inst_cell_102_49 ( BL49, BLN49, WL102);
sram_cell_6t_3 inst_cell_102_48 ( BL48, BLN48, WL102);
sram_cell_6t_3 inst_cell_102_47 ( BL47, BLN47, WL102);
sram_cell_6t_3 inst_cell_102_46 ( BL46, BLN46, WL102);
sram_cell_6t_3 inst_cell_102_45 ( BL45, BLN45, WL102);
sram_cell_6t_3 inst_cell_102_44 ( BL44, BLN44, WL102);
sram_cell_6t_3 inst_cell_102_43 ( BL43, BLN43, WL102);
sram_cell_6t_3 inst_cell_102_42 ( BL42, BLN42, WL102);
sram_cell_6t_3 inst_cell_102_41 ( BL41, BLN41, WL102);
sram_cell_6t_3 inst_cell_102_40 ( BL40, BLN40, WL102);
sram_cell_6t_3 inst_cell_102_39 ( BL39, BLN39, WL102);
sram_cell_6t_3 inst_cell_102_38 ( BL38, BLN38, WL102);
sram_cell_6t_3 inst_cell_102_37 ( BL37, BLN37, WL102);
sram_cell_6t_3 inst_cell_102_36 ( BL36, BLN36, WL102);
sram_cell_6t_3 inst_cell_102_35 ( BL35, BLN35, WL102);
sram_cell_6t_3 inst_cell_102_34 ( BL34, BLN34, WL102);
sram_cell_6t_3 inst_cell_102_33 ( BL33, BLN33, WL102);
sram_cell_6t_3 inst_cell_102_32 ( BL32, BLN32, WL102);
sram_cell_6t_3 inst_cell_102_31 ( BL31, BLN31, WL102);
sram_cell_6t_3 inst_cell_102_30 ( BL30, BLN30, WL102);
sram_cell_6t_3 inst_cell_102_29 ( BL29, BLN29, WL102);
sram_cell_6t_3 inst_cell_102_28 ( BL28, BLN28, WL102);
sram_cell_6t_3 inst_cell_102_27 ( BL27, BLN27, WL102);
sram_cell_6t_3 inst_cell_102_26 ( BL26, BLN26, WL102);
sram_cell_6t_3 inst_cell_102_25 ( BL25, BLN25, WL102);
sram_cell_6t_3 inst_cell_102_24 ( BL24, BLN24, WL102);
sram_cell_6t_3 inst_cell_102_23 ( BL23, BLN23, WL102);
sram_cell_6t_3 inst_cell_102_22 ( BL22, BLN22, WL102);
sram_cell_6t_3 inst_cell_102_21 ( BL21, BLN21, WL102);
sram_cell_6t_3 inst_cell_102_20 ( BL20, BLN20, WL102);
sram_cell_6t_3 inst_cell_102_19 ( BL19, BLN19, WL102);
sram_cell_6t_3 inst_cell_102_18 ( BL18, BLN18, WL102);
sram_cell_6t_3 inst_cell_102_17 ( BL17, BLN17, WL102);
sram_cell_6t_3 inst_cell_102_16 ( BL16, BLN16, WL102);
sram_cell_6t_3 inst_cell_102_15 ( BL15, BLN15, WL102);
sram_cell_6t_3 inst_cell_102_14 ( BL14, BLN14, WL102);
sram_cell_6t_3 inst_cell_102_13 ( BL13, BLN13, WL102);
sram_cell_6t_3 inst_cell_102_12 ( BL12, BLN12, WL102);
sram_cell_6t_3 inst_cell_102_11 ( BL11, BLN11, WL102);
sram_cell_6t_3 inst_cell_102_10 ( BL10, BLN10, WL102);
sram_cell_6t_3 inst_cell_102_9 ( BL9, BLN9, WL102);
sram_cell_6t_3 inst_cell_102_8 ( BL8, BLN8, WL102);
sram_cell_6t_3 inst_cell_102_7 ( BL7, BLN7, WL102);
sram_cell_6t_3 inst_cell_102_6 ( BL6, BLN6, WL102);
sram_cell_6t_3 inst_cell_102_5 ( BL5, BLN5, WL102);
sram_cell_6t_3 inst_cell_102_4 ( BL4, BLN4, WL102);
sram_cell_6t_3 inst_cell_102_3 ( BL3, BLN3, WL102);
sram_cell_6t_3 inst_cell_102_2 ( BL2, BLN2, WL102);
sram_cell_6t_3 inst_cell_102_1 ( BL1, BLN1, WL102);
sram_cell_6t_3 inst_cell_102_0 ( BL0, BLN0, WL102);
sram_cell_6t_3 inst_cell_101_127 ( BL127, BLN127, WL101);
sram_cell_6t_3 inst_cell_101_126 ( BL126, BLN126, WL101);
sram_cell_6t_3 inst_cell_101_125 ( BL125, BLN125, WL101);
sram_cell_6t_3 inst_cell_101_124 ( BL124, BLN124, WL101);
sram_cell_6t_3 inst_cell_101_123 ( BL123, BLN123, WL101);
sram_cell_6t_3 inst_cell_101_122 ( BL122, BLN122, WL101);
sram_cell_6t_3 inst_cell_101_121 ( BL121, BLN121, WL101);
sram_cell_6t_3 inst_cell_101_120 ( BL120, BLN120, WL101);
sram_cell_6t_3 inst_cell_101_119 ( BL119, BLN119, WL101);
sram_cell_6t_3 inst_cell_101_118 ( BL118, BLN118, WL101);
sram_cell_6t_3 inst_cell_101_117 ( BL117, BLN117, WL101);
sram_cell_6t_3 inst_cell_101_116 ( BL116, BLN116, WL101);
sram_cell_6t_3 inst_cell_101_115 ( BL115, BLN115, WL101);
sram_cell_6t_3 inst_cell_101_114 ( BL114, BLN114, WL101);
sram_cell_6t_3 inst_cell_101_113 ( BL113, BLN113, WL101);
sram_cell_6t_3 inst_cell_101_112 ( BL112, BLN112, WL101);
sram_cell_6t_3 inst_cell_101_111 ( BL111, BLN111, WL101);
sram_cell_6t_3 inst_cell_101_110 ( BL110, BLN110, WL101);
sram_cell_6t_3 inst_cell_101_109 ( BL109, BLN109, WL101);
sram_cell_6t_3 inst_cell_101_108 ( BL108, BLN108, WL101);
sram_cell_6t_3 inst_cell_101_107 ( BL107, BLN107, WL101);
sram_cell_6t_3 inst_cell_101_106 ( BL106, BLN106, WL101);
sram_cell_6t_3 inst_cell_101_105 ( BL105, BLN105, WL101);
sram_cell_6t_3 inst_cell_101_104 ( BL104, BLN104, WL101);
sram_cell_6t_3 inst_cell_101_103 ( BL103, BLN103, WL101);
sram_cell_6t_3 inst_cell_101_102 ( BL102, BLN102, WL101);
sram_cell_6t_3 inst_cell_101_101 ( BL101, BLN101, WL101);
sram_cell_6t_3 inst_cell_101_100 ( BL100, BLN100, WL101);
sram_cell_6t_3 inst_cell_101_99 ( BL99, BLN99, WL101);
sram_cell_6t_3 inst_cell_101_98 ( BL98, BLN98, WL101);
sram_cell_6t_3 inst_cell_101_97 ( BL97, BLN97, WL101);
sram_cell_6t_3 inst_cell_101_96 ( BL96, BLN96, WL101);
sram_cell_6t_3 inst_cell_101_95 ( BL95, BLN95, WL101);
sram_cell_6t_3 inst_cell_101_94 ( BL94, BLN94, WL101);
sram_cell_6t_3 inst_cell_101_93 ( BL93, BLN93, WL101);
sram_cell_6t_3 inst_cell_101_92 ( BL92, BLN92, WL101);
sram_cell_6t_3 inst_cell_101_91 ( BL91, BLN91, WL101);
sram_cell_6t_3 inst_cell_101_90 ( BL90, BLN90, WL101);
sram_cell_6t_3 inst_cell_101_89 ( BL89, BLN89, WL101);
sram_cell_6t_3 inst_cell_101_88 ( BL88, BLN88, WL101);
sram_cell_6t_3 inst_cell_101_87 ( BL87, BLN87, WL101);
sram_cell_6t_3 inst_cell_101_86 ( BL86, BLN86, WL101);
sram_cell_6t_3 inst_cell_101_85 ( BL85, BLN85, WL101);
sram_cell_6t_3 inst_cell_101_84 ( BL84, BLN84, WL101);
sram_cell_6t_3 inst_cell_101_83 ( BL83, BLN83, WL101);
sram_cell_6t_3 inst_cell_101_82 ( BL82, BLN82, WL101);
sram_cell_6t_3 inst_cell_101_81 ( BL81, BLN81, WL101);
sram_cell_6t_3 inst_cell_101_80 ( BL80, BLN80, WL101);
sram_cell_6t_3 inst_cell_101_79 ( BL79, BLN79, WL101);
sram_cell_6t_3 inst_cell_101_78 ( BL78, BLN78, WL101);
sram_cell_6t_3 inst_cell_101_77 ( BL77, BLN77, WL101);
sram_cell_6t_3 inst_cell_101_76 ( BL76, BLN76, WL101);
sram_cell_6t_3 inst_cell_101_75 ( BL75, BLN75, WL101);
sram_cell_6t_3 inst_cell_101_74 ( BL74, BLN74, WL101);
sram_cell_6t_3 inst_cell_101_73 ( BL73, BLN73, WL101);
sram_cell_6t_3 inst_cell_101_72 ( BL72, BLN72, WL101);
sram_cell_6t_3 inst_cell_101_71 ( BL71, BLN71, WL101);
sram_cell_6t_3 inst_cell_101_70 ( BL70, BLN70, WL101);
sram_cell_6t_3 inst_cell_101_69 ( BL69, BLN69, WL101);
sram_cell_6t_3 inst_cell_101_68 ( BL68, BLN68, WL101);
sram_cell_6t_3 inst_cell_101_67 ( BL67, BLN67, WL101);
sram_cell_6t_3 inst_cell_101_66 ( BL66, BLN66, WL101);
sram_cell_6t_3 inst_cell_101_65 ( BL65, BLN65, WL101);
sram_cell_6t_3 inst_cell_101_64 ( BL64, BLN64, WL101);
sram_cell_6t_3 inst_cell_101_63 ( BL63, BLN63, WL101);
sram_cell_6t_3 inst_cell_101_62 ( BL62, BLN62, WL101);
sram_cell_6t_3 inst_cell_101_61 ( BL61, BLN61, WL101);
sram_cell_6t_3 inst_cell_101_60 ( BL60, BLN60, WL101);
sram_cell_6t_3 inst_cell_101_59 ( BL59, BLN59, WL101);
sram_cell_6t_3 inst_cell_101_58 ( BL58, BLN58, WL101);
sram_cell_6t_3 inst_cell_101_57 ( BL57, BLN57, WL101);
sram_cell_6t_3 inst_cell_101_56 ( BL56, BLN56, WL101);
sram_cell_6t_3 inst_cell_101_55 ( BL55, BLN55, WL101);
sram_cell_6t_3 inst_cell_101_54 ( BL54, BLN54, WL101);
sram_cell_6t_3 inst_cell_101_53 ( BL53, BLN53, WL101);
sram_cell_6t_3 inst_cell_101_52 ( BL52, BLN52, WL101);
sram_cell_6t_3 inst_cell_101_51 ( BL51, BLN51, WL101);
sram_cell_6t_3 inst_cell_101_50 ( BL50, BLN50, WL101);
sram_cell_6t_3 inst_cell_101_49 ( BL49, BLN49, WL101);
sram_cell_6t_3 inst_cell_101_48 ( BL48, BLN48, WL101);
sram_cell_6t_3 inst_cell_101_47 ( BL47, BLN47, WL101);
sram_cell_6t_3 inst_cell_101_46 ( BL46, BLN46, WL101);
sram_cell_6t_3 inst_cell_101_45 ( BL45, BLN45, WL101);
sram_cell_6t_3 inst_cell_101_44 ( BL44, BLN44, WL101);
sram_cell_6t_3 inst_cell_101_43 ( BL43, BLN43, WL101);
sram_cell_6t_3 inst_cell_101_42 ( BL42, BLN42, WL101);
sram_cell_6t_3 inst_cell_101_41 ( BL41, BLN41, WL101);
sram_cell_6t_3 inst_cell_101_40 ( BL40, BLN40, WL101);
sram_cell_6t_3 inst_cell_101_39 ( BL39, BLN39, WL101);
sram_cell_6t_3 inst_cell_101_38 ( BL38, BLN38, WL101);
sram_cell_6t_3 inst_cell_101_37 ( BL37, BLN37, WL101);
sram_cell_6t_3 inst_cell_101_36 ( BL36, BLN36, WL101);
sram_cell_6t_3 inst_cell_101_35 ( BL35, BLN35, WL101);
sram_cell_6t_3 inst_cell_101_34 ( BL34, BLN34, WL101);
sram_cell_6t_3 inst_cell_101_33 ( BL33, BLN33, WL101);
sram_cell_6t_3 inst_cell_101_32 ( BL32, BLN32, WL101);
sram_cell_6t_3 inst_cell_101_31 ( BL31, BLN31, WL101);
sram_cell_6t_3 inst_cell_101_30 ( BL30, BLN30, WL101);
sram_cell_6t_3 inst_cell_101_29 ( BL29, BLN29, WL101);
sram_cell_6t_3 inst_cell_101_28 ( BL28, BLN28, WL101);
sram_cell_6t_3 inst_cell_101_27 ( BL27, BLN27, WL101);
sram_cell_6t_3 inst_cell_101_26 ( BL26, BLN26, WL101);
sram_cell_6t_3 inst_cell_101_25 ( BL25, BLN25, WL101);
sram_cell_6t_3 inst_cell_101_24 ( BL24, BLN24, WL101);
sram_cell_6t_3 inst_cell_101_23 ( BL23, BLN23, WL101);
sram_cell_6t_3 inst_cell_101_22 ( BL22, BLN22, WL101);
sram_cell_6t_3 inst_cell_101_21 ( BL21, BLN21, WL101);
sram_cell_6t_3 inst_cell_101_20 ( BL20, BLN20, WL101);
sram_cell_6t_3 inst_cell_101_19 ( BL19, BLN19, WL101);
sram_cell_6t_3 inst_cell_101_18 ( BL18, BLN18, WL101);
sram_cell_6t_3 inst_cell_101_17 ( BL17, BLN17, WL101);
sram_cell_6t_3 inst_cell_101_16 ( BL16, BLN16, WL101);
sram_cell_6t_3 inst_cell_101_15 ( BL15, BLN15, WL101);
sram_cell_6t_3 inst_cell_101_14 ( BL14, BLN14, WL101);
sram_cell_6t_3 inst_cell_101_13 ( BL13, BLN13, WL101);
sram_cell_6t_3 inst_cell_101_12 ( BL12, BLN12, WL101);
sram_cell_6t_3 inst_cell_101_11 ( BL11, BLN11, WL101);
sram_cell_6t_3 inst_cell_101_10 ( BL10, BLN10, WL101);
sram_cell_6t_3 inst_cell_101_9 ( BL9, BLN9, WL101);
sram_cell_6t_3 inst_cell_101_8 ( BL8, BLN8, WL101);
sram_cell_6t_3 inst_cell_101_7 ( BL7, BLN7, WL101);
sram_cell_6t_3 inst_cell_101_6 ( BL6, BLN6, WL101);
sram_cell_6t_3 inst_cell_101_5 ( BL5, BLN5, WL101);
sram_cell_6t_3 inst_cell_101_4 ( BL4, BLN4, WL101);
sram_cell_6t_3 inst_cell_101_3 ( BL3, BLN3, WL101);
sram_cell_6t_3 inst_cell_101_2 ( BL2, BLN2, WL101);
sram_cell_6t_3 inst_cell_101_1 ( BL1, BLN1, WL101);
sram_cell_6t_3 inst_cell_101_0 ( BL0, BLN0, WL101);
sram_cell_6t_3 inst_cell_100_127 ( BL127, BLN127, WL100);
sram_cell_6t_3 inst_cell_100_126 ( BL126, BLN126, WL100);
sram_cell_6t_3 inst_cell_100_125 ( BL125, BLN125, WL100);
sram_cell_6t_3 inst_cell_100_124 ( BL124, BLN124, WL100);
sram_cell_6t_3 inst_cell_100_123 ( BL123, BLN123, WL100);
sram_cell_6t_3 inst_cell_100_122 ( BL122, BLN122, WL100);
sram_cell_6t_3 inst_cell_100_121 ( BL121, BLN121, WL100);
sram_cell_6t_3 inst_cell_100_120 ( BL120, BLN120, WL100);
sram_cell_6t_3 inst_cell_100_119 ( BL119, BLN119, WL100);
sram_cell_6t_3 inst_cell_100_118 ( BL118, BLN118, WL100);
sram_cell_6t_3 inst_cell_100_117 ( BL117, BLN117, WL100);
sram_cell_6t_3 inst_cell_100_116 ( BL116, BLN116, WL100);
sram_cell_6t_3 inst_cell_100_115 ( BL115, BLN115, WL100);
sram_cell_6t_3 inst_cell_100_114 ( BL114, BLN114, WL100);
sram_cell_6t_3 inst_cell_100_113 ( BL113, BLN113, WL100);
sram_cell_6t_3 inst_cell_100_112 ( BL112, BLN112, WL100);
sram_cell_6t_3 inst_cell_100_111 ( BL111, BLN111, WL100);
sram_cell_6t_3 inst_cell_100_110 ( BL110, BLN110, WL100);
sram_cell_6t_3 inst_cell_100_109 ( BL109, BLN109, WL100);
sram_cell_6t_3 inst_cell_100_108 ( BL108, BLN108, WL100);
sram_cell_6t_3 inst_cell_100_107 ( BL107, BLN107, WL100);
sram_cell_6t_3 inst_cell_100_106 ( BL106, BLN106, WL100);
sram_cell_6t_3 inst_cell_100_105 ( BL105, BLN105, WL100);
sram_cell_6t_3 inst_cell_100_104 ( BL104, BLN104, WL100);
sram_cell_6t_3 inst_cell_100_103 ( BL103, BLN103, WL100);
sram_cell_6t_3 inst_cell_100_102 ( BL102, BLN102, WL100);
sram_cell_6t_3 inst_cell_100_101 ( BL101, BLN101, WL100);
sram_cell_6t_3 inst_cell_100_100 ( BL100, BLN100, WL100);
sram_cell_6t_3 inst_cell_100_99 ( BL99, BLN99, WL100);
sram_cell_6t_3 inst_cell_100_98 ( BL98, BLN98, WL100);
sram_cell_6t_3 inst_cell_100_97 ( BL97, BLN97, WL100);
sram_cell_6t_3 inst_cell_100_96 ( BL96, BLN96, WL100);
sram_cell_6t_3 inst_cell_100_95 ( BL95, BLN95, WL100);
sram_cell_6t_3 inst_cell_100_94 ( BL94, BLN94, WL100);
sram_cell_6t_3 inst_cell_100_93 ( BL93, BLN93, WL100);
sram_cell_6t_3 inst_cell_100_92 ( BL92, BLN92, WL100);
sram_cell_6t_3 inst_cell_100_91 ( BL91, BLN91, WL100);
sram_cell_6t_3 inst_cell_100_90 ( BL90, BLN90, WL100);
sram_cell_6t_3 inst_cell_100_89 ( BL89, BLN89, WL100);
sram_cell_6t_3 inst_cell_100_88 ( BL88, BLN88, WL100);
sram_cell_6t_3 inst_cell_100_87 ( BL87, BLN87, WL100);
sram_cell_6t_3 inst_cell_100_86 ( BL86, BLN86, WL100);
sram_cell_6t_3 inst_cell_100_85 ( BL85, BLN85, WL100);
sram_cell_6t_3 inst_cell_100_84 ( BL84, BLN84, WL100);
sram_cell_6t_3 inst_cell_100_83 ( BL83, BLN83, WL100);
sram_cell_6t_3 inst_cell_100_82 ( BL82, BLN82, WL100);
sram_cell_6t_3 inst_cell_100_81 ( BL81, BLN81, WL100);
sram_cell_6t_3 inst_cell_100_80 ( BL80, BLN80, WL100);
sram_cell_6t_3 inst_cell_100_79 ( BL79, BLN79, WL100);
sram_cell_6t_3 inst_cell_100_78 ( BL78, BLN78, WL100);
sram_cell_6t_3 inst_cell_100_77 ( BL77, BLN77, WL100);
sram_cell_6t_3 inst_cell_100_76 ( BL76, BLN76, WL100);
sram_cell_6t_3 inst_cell_100_75 ( BL75, BLN75, WL100);
sram_cell_6t_3 inst_cell_100_74 ( BL74, BLN74, WL100);
sram_cell_6t_3 inst_cell_100_73 ( BL73, BLN73, WL100);
sram_cell_6t_3 inst_cell_100_72 ( BL72, BLN72, WL100);
sram_cell_6t_3 inst_cell_100_71 ( BL71, BLN71, WL100);
sram_cell_6t_3 inst_cell_100_70 ( BL70, BLN70, WL100);
sram_cell_6t_3 inst_cell_100_69 ( BL69, BLN69, WL100);
sram_cell_6t_3 inst_cell_100_68 ( BL68, BLN68, WL100);
sram_cell_6t_3 inst_cell_100_67 ( BL67, BLN67, WL100);
sram_cell_6t_3 inst_cell_100_66 ( BL66, BLN66, WL100);
sram_cell_6t_3 inst_cell_100_65 ( BL65, BLN65, WL100);
sram_cell_6t_3 inst_cell_100_64 ( BL64, BLN64, WL100);
sram_cell_6t_3 inst_cell_100_63 ( BL63, BLN63, WL100);
sram_cell_6t_3 inst_cell_100_62 ( BL62, BLN62, WL100);
sram_cell_6t_3 inst_cell_100_61 ( BL61, BLN61, WL100);
sram_cell_6t_3 inst_cell_100_60 ( BL60, BLN60, WL100);
sram_cell_6t_3 inst_cell_100_59 ( BL59, BLN59, WL100);
sram_cell_6t_3 inst_cell_100_58 ( BL58, BLN58, WL100);
sram_cell_6t_3 inst_cell_100_57 ( BL57, BLN57, WL100);
sram_cell_6t_3 inst_cell_100_56 ( BL56, BLN56, WL100);
sram_cell_6t_3 inst_cell_100_55 ( BL55, BLN55, WL100);
sram_cell_6t_3 inst_cell_100_54 ( BL54, BLN54, WL100);
sram_cell_6t_3 inst_cell_100_53 ( BL53, BLN53, WL100);
sram_cell_6t_3 inst_cell_100_52 ( BL52, BLN52, WL100);
sram_cell_6t_3 inst_cell_100_51 ( BL51, BLN51, WL100);
sram_cell_6t_3 inst_cell_100_50 ( BL50, BLN50, WL100);
sram_cell_6t_3 inst_cell_100_49 ( BL49, BLN49, WL100);
sram_cell_6t_3 inst_cell_100_48 ( BL48, BLN48, WL100);
sram_cell_6t_3 inst_cell_100_47 ( BL47, BLN47, WL100);
sram_cell_6t_3 inst_cell_100_46 ( BL46, BLN46, WL100);
sram_cell_6t_3 inst_cell_100_45 ( BL45, BLN45, WL100);
sram_cell_6t_3 inst_cell_100_44 ( BL44, BLN44, WL100);
sram_cell_6t_3 inst_cell_100_43 ( BL43, BLN43, WL100);
sram_cell_6t_3 inst_cell_100_42 ( BL42, BLN42, WL100);
sram_cell_6t_3 inst_cell_100_41 ( BL41, BLN41, WL100);
sram_cell_6t_3 inst_cell_100_40 ( BL40, BLN40, WL100);
sram_cell_6t_3 inst_cell_100_39 ( BL39, BLN39, WL100);
sram_cell_6t_3 inst_cell_100_38 ( BL38, BLN38, WL100);
sram_cell_6t_3 inst_cell_100_37 ( BL37, BLN37, WL100);
sram_cell_6t_3 inst_cell_100_36 ( BL36, BLN36, WL100);
sram_cell_6t_3 inst_cell_100_35 ( BL35, BLN35, WL100);
sram_cell_6t_3 inst_cell_100_34 ( BL34, BLN34, WL100);
sram_cell_6t_3 inst_cell_100_33 ( BL33, BLN33, WL100);
sram_cell_6t_3 inst_cell_100_32 ( BL32, BLN32, WL100);
sram_cell_6t_3 inst_cell_100_31 ( BL31, BLN31, WL100);
sram_cell_6t_3 inst_cell_100_30 ( BL30, BLN30, WL100);
sram_cell_6t_3 inst_cell_100_29 ( BL29, BLN29, WL100);
sram_cell_6t_3 inst_cell_100_28 ( BL28, BLN28, WL100);
sram_cell_6t_3 inst_cell_100_27 ( BL27, BLN27, WL100);
sram_cell_6t_3 inst_cell_100_26 ( BL26, BLN26, WL100);
sram_cell_6t_3 inst_cell_100_25 ( BL25, BLN25, WL100);
sram_cell_6t_3 inst_cell_100_24 ( BL24, BLN24, WL100);
sram_cell_6t_3 inst_cell_100_23 ( BL23, BLN23, WL100);
sram_cell_6t_3 inst_cell_100_22 ( BL22, BLN22, WL100);
sram_cell_6t_3 inst_cell_100_21 ( BL21, BLN21, WL100);
sram_cell_6t_3 inst_cell_100_20 ( BL20, BLN20, WL100);
sram_cell_6t_3 inst_cell_100_19 ( BL19, BLN19, WL100);
sram_cell_6t_3 inst_cell_100_18 ( BL18, BLN18, WL100);
sram_cell_6t_3 inst_cell_100_17 ( BL17, BLN17, WL100);
sram_cell_6t_3 inst_cell_100_16 ( BL16, BLN16, WL100);
sram_cell_6t_3 inst_cell_100_15 ( BL15, BLN15, WL100);
sram_cell_6t_3 inst_cell_100_14 ( BL14, BLN14, WL100);
sram_cell_6t_3 inst_cell_100_13 ( BL13, BLN13, WL100);
sram_cell_6t_3 inst_cell_100_12 ( BL12, BLN12, WL100);
sram_cell_6t_3 inst_cell_100_11 ( BL11, BLN11, WL100);
sram_cell_6t_3 inst_cell_100_10 ( BL10, BLN10, WL100);
sram_cell_6t_3 inst_cell_100_9 ( BL9, BLN9, WL100);
sram_cell_6t_3 inst_cell_100_8 ( BL8, BLN8, WL100);
sram_cell_6t_3 inst_cell_100_7 ( BL7, BLN7, WL100);
sram_cell_6t_3 inst_cell_100_6 ( BL6, BLN6, WL100);
sram_cell_6t_3 inst_cell_100_5 ( BL5, BLN5, WL100);
sram_cell_6t_3 inst_cell_100_4 ( BL4, BLN4, WL100);
sram_cell_6t_3 inst_cell_100_3 ( BL3, BLN3, WL100);
sram_cell_6t_3 inst_cell_100_2 ( BL2, BLN2, WL100);
sram_cell_6t_3 inst_cell_100_1 ( BL1, BLN1, WL100);
sram_cell_6t_3 inst_cell_100_0 ( BL0, BLN0, WL100);
sram_cell_6t_3 inst_cell_99_127 ( BL127, BLN127, WL99);
sram_cell_6t_3 inst_cell_99_126 ( BL126, BLN126, WL99);
sram_cell_6t_3 inst_cell_99_125 ( BL125, BLN125, WL99);
sram_cell_6t_3 inst_cell_99_124 ( BL124, BLN124, WL99);
sram_cell_6t_3 inst_cell_99_123 ( BL123, BLN123, WL99);
sram_cell_6t_3 inst_cell_99_122 ( BL122, BLN122, WL99);
sram_cell_6t_3 inst_cell_99_121 ( BL121, BLN121, WL99);
sram_cell_6t_3 inst_cell_99_120 ( BL120, BLN120, WL99);
sram_cell_6t_3 inst_cell_99_119 ( BL119, BLN119, WL99);
sram_cell_6t_3 inst_cell_99_118 ( BL118, BLN118, WL99);
sram_cell_6t_3 inst_cell_99_117 ( BL117, BLN117, WL99);
sram_cell_6t_3 inst_cell_99_116 ( BL116, BLN116, WL99);
sram_cell_6t_3 inst_cell_99_115 ( BL115, BLN115, WL99);
sram_cell_6t_3 inst_cell_99_114 ( BL114, BLN114, WL99);
sram_cell_6t_3 inst_cell_99_113 ( BL113, BLN113, WL99);
sram_cell_6t_3 inst_cell_99_112 ( BL112, BLN112, WL99);
sram_cell_6t_3 inst_cell_99_111 ( BL111, BLN111, WL99);
sram_cell_6t_3 inst_cell_99_110 ( BL110, BLN110, WL99);
sram_cell_6t_3 inst_cell_99_109 ( BL109, BLN109, WL99);
sram_cell_6t_3 inst_cell_99_108 ( BL108, BLN108, WL99);
sram_cell_6t_3 inst_cell_99_107 ( BL107, BLN107, WL99);
sram_cell_6t_3 inst_cell_99_106 ( BL106, BLN106, WL99);
sram_cell_6t_3 inst_cell_99_105 ( BL105, BLN105, WL99);
sram_cell_6t_3 inst_cell_99_104 ( BL104, BLN104, WL99);
sram_cell_6t_3 inst_cell_99_103 ( BL103, BLN103, WL99);
sram_cell_6t_3 inst_cell_99_102 ( BL102, BLN102, WL99);
sram_cell_6t_3 inst_cell_99_101 ( BL101, BLN101, WL99);
sram_cell_6t_3 inst_cell_99_100 ( BL100, BLN100, WL99);
sram_cell_6t_3 inst_cell_99_99 ( BL99, BLN99, WL99);
sram_cell_6t_3 inst_cell_99_98 ( BL98, BLN98, WL99);
sram_cell_6t_3 inst_cell_99_97 ( BL97, BLN97, WL99);
sram_cell_6t_3 inst_cell_99_96 ( BL96, BLN96, WL99);
sram_cell_6t_3 inst_cell_99_95 ( BL95, BLN95, WL99);
sram_cell_6t_3 inst_cell_99_94 ( BL94, BLN94, WL99);
sram_cell_6t_3 inst_cell_99_93 ( BL93, BLN93, WL99);
sram_cell_6t_3 inst_cell_99_92 ( BL92, BLN92, WL99);
sram_cell_6t_3 inst_cell_99_91 ( BL91, BLN91, WL99);
sram_cell_6t_3 inst_cell_99_90 ( BL90, BLN90, WL99);
sram_cell_6t_3 inst_cell_99_89 ( BL89, BLN89, WL99);
sram_cell_6t_3 inst_cell_99_88 ( BL88, BLN88, WL99);
sram_cell_6t_3 inst_cell_99_87 ( BL87, BLN87, WL99);
sram_cell_6t_3 inst_cell_99_86 ( BL86, BLN86, WL99);
sram_cell_6t_3 inst_cell_99_85 ( BL85, BLN85, WL99);
sram_cell_6t_3 inst_cell_99_84 ( BL84, BLN84, WL99);
sram_cell_6t_3 inst_cell_99_83 ( BL83, BLN83, WL99);
sram_cell_6t_3 inst_cell_99_82 ( BL82, BLN82, WL99);
sram_cell_6t_3 inst_cell_99_81 ( BL81, BLN81, WL99);
sram_cell_6t_3 inst_cell_99_80 ( BL80, BLN80, WL99);
sram_cell_6t_3 inst_cell_99_79 ( BL79, BLN79, WL99);
sram_cell_6t_3 inst_cell_99_78 ( BL78, BLN78, WL99);
sram_cell_6t_3 inst_cell_99_77 ( BL77, BLN77, WL99);
sram_cell_6t_3 inst_cell_99_76 ( BL76, BLN76, WL99);
sram_cell_6t_3 inst_cell_99_75 ( BL75, BLN75, WL99);
sram_cell_6t_3 inst_cell_99_74 ( BL74, BLN74, WL99);
sram_cell_6t_3 inst_cell_99_73 ( BL73, BLN73, WL99);
sram_cell_6t_3 inst_cell_99_72 ( BL72, BLN72, WL99);
sram_cell_6t_3 inst_cell_99_71 ( BL71, BLN71, WL99);
sram_cell_6t_3 inst_cell_99_70 ( BL70, BLN70, WL99);
sram_cell_6t_3 inst_cell_99_69 ( BL69, BLN69, WL99);
sram_cell_6t_3 inst_cell_99_68 ( BL68, BLN68, WL99);
sram_cell_6t_3 inst_cell_99_67 ( BL67, BLN67, WL99);
sram_cell_6t_3 inst_cell_99_66 ( BL66, BLN66, WL99);
sram_cell_6t_3 inst_cell_99_65 ( BL65, BLN65, WL99);
sram_cell_6t_3 inst_cell_99_64 ( BL64, BLN64, WL99);
sram_cell_6t_3 inst_cell_99_63 ( BL63, BLN63, WL99);
sram_cell_6t_3 inst_cell_99_62 ( BL62, BLN62, WL99);
sram_cell_6t_3 inst_cell_99_61 ( BL61, BLN61, WL99);
sram_cell_6t_3 inst_cell_99_60 ( BL60, BLN60, WL99);
sram_cell_6t_3 inst_cell_99_59 ( BL59, BLN59, WL99);
sram_cell_6t_3 inst_cell_99_58 ( BL58, BLN58, WL99);
sram_cell_6t_3 inst_cell_99_57 ( BL57, BLN57, WL99);
sram_cell_6t_3 inst_cell_99_56 ( BL56, BLN56, WL99);
sram_cell_6t_3 inst_cell_99_55 ( BL55, BLN55, WL99);
sram_cell_6t_3 inst_cell_99_54 ( BL54, BLN54, WL99);
sram_cell_6t_3 inst_cell_99_53 ( BL53, BLN53, WL99);
sram_cell_6t_3 inst_cell_99_52 ( BL52, BLN52, WL99);
sram_cell_6t_3 inst_cell_99_51 ( BL51, BLN51, WL99);
sram_cell_6t_3 inst_cell_99_50 ( BL50, BLN50, WL99);
sram_cell_6t_3 inst_cell_99_49 ( BL49, BLN49, WL99);
sram_cell_6t_3 inst_cell_99_48 ( BL48, BLN48, WL99);
sram_cell_6t_3 inst_cell_99_47 ( BL47, BLN47, WL99);
sram_cell_6t_3 inst_cell_99_46 ( BL46, BLN46, WL99);
sram_cell_6t_3 inst_cell_99_45 ( BL45, BLN45, WL99);
sram_cell_6t_3 inst_cell_99_44 ( BL44, BLN44, WL99);
sram_cell_6t_3 inst_cell_99_43 ( BL43, BLN43, WL99);
sram_cell_6t_3 inst_cell_99_42 ( BL42, BLN42, WL99);
sram_cell_6t_3 inst_cell_99_41 ( BL41, BLN41, WL99);
sram_cell_6t_3 inst_cell_99_40 ( BL40, BLN40, WL99);
sram_cell_6t_3 inst_cell_99_39 ( BL39, BLN39, WL99);
sram_cell_6t_3 inst_cell_99_38 ( BL38, BLN38, WL99);
sram_cell_6t_3 inst_cell_99_37 ( BL37, BLN37, WL99);
sram_cell_6t_3 inst_cell_99_36 ( BL36, BLN36, WL99);
sram_cell_6t_3 inst_cell_99_35 ( BL35, BLN35, WL99);
sram_cell_6t_3 inst_cell_99_34 ( BL34, BLN34, WL99);
sram_cell_6t_3 inst_cell_99_33 ( BL33, BLN33, WL99);
sram_cell_6t_3 inst_cell_99_32 ( BL32, BLN32, WL99);
sram_cell_6t_3 inst_cell_99_31 ( BL31, BLN31, WL99);
sram_cell_6t_3 inst_cell_99_30 ( BL30, BLN30, WL99);
sram_cell_6t_3 inst_cell_99_29 ( BL29, BLN29, WL99);
sram_cell_6t_3 inst_cell_99_28 ( BL28, BLN28, WL99);
sram_cell_6t_3 inst_cell_99_27 ( BL27, BLN27, WL99);
sram_cell_6t_3 inst_cell_99_26 ( BL26, BLN26, WL99);
sram_cell_6t_3 inst_cell_99_25 ( BL25, BLN25, WL99);
sram_cell_6t_3 inst_cell_99_24 ( BL24, BLN24, WL99);
sram_cell_6t_3 inst_cell_99_23 ( BL23, BLN23, WL99);
sram_cell_6t_3 inst_cell_99_22 ( BL22, BLN22, WL99);
sram_cell_6t_3 inst_cell_99_21 ( BL21, BLN21, WL99);
sram_cell_6t_3 inst_cell_99_20 ( BL20, BLN20, WL99);
sram_cell_6t_3 inst_cell_99_19 ( BL19, BLN19, WL99);
sram_cell_6t_3 inst_cell_99_18 ( BL18, BLN18, WL99);
sram_cell_6t_3 inst_cell_99_17 ( BL17, BLN17, WL99);
sram_cell_6t_3 inst_cell_99_16 ( BL16, BLN16, WL99);
sram_cell_6t_3 inst_cell_99_15 ( BL15, BLN15, WL99);
sram_cell_6t_3 inst_cell_99_14 ( BL14, BLN14, WL99);
sram_cell_6t_3 inst_cell_99_13 ( BL13, BLN13, WL99);
sram_cell_6t_3 inst_cell_99_12 ( BL12, BLN12, WL99);
sram_cell_6t_3 inst_cell_99_11 ( BL11, BLN11, WL99);
sram_cell_6t_3 inst_cell_99_10 ( BL10, BLN10, WL99);
sram_cell_6t_3 inst_cell_99_9 ( BL9, BLN9, WL99);
sram_cell_6t_3 inst_cell_99_8 ( BL8, BLN8, WL99);
sram_cell_6t_3 inst_cell_99_7 ( BL7, BLN7, WL99);
sram_cell_6t_3 inst_cell_99_6 ( BL6, BLN6, WL99);
sram_cell_6t_3 inst_cell_99_5 ( BL5, BLN5, WL99);
sram_cell_6t_3 inst_cell_99_4 ( BL4, BLN4, WL99);
sram_cell_6t_3 inst_cell_99_3 ( BL3, BLN3, WL99);
sram_cell_6t_3 inst_cell_99_2 ( BL2, BLN2, WL99);
sram_cell_6t_3 inst_cell_99_1 ( BL1, BLN1, WL99);
sram_cell_6t_3 inst_cell_99_0 ( BL0, BLN0, WL99);
sram_cell_6t_3 inst_cell_98_127 ( BL127, BLN127, WL98);
sram_cell_6t_3 inst_cell_98_126 ( BL126, BLN126, WL98);
sram_cell_6t_3 inst_cell_98_125 ( BL125, BLN125, WL98);
sram_cell_6t_3 inst_cell_98_124 ( BL124, BLN124, WL98);
sram_cell_6t_3 inst_cell_98_123 ( BL123, BLN123, WL98);
sram_cell_6t_3 inst_cell_98_122 ( BL122, BLN122, WL98);
sram_cell_6t_3 inst_cell_98_121 ( BL121, BLN121, WL98);
sram_cell_6t_3 inst_cell_98_120 ( BL120, BLN120, WL98);
sram_cell_6t_3 inst_cell_98_119 ( BL119, BLN119, WL98);
sram_cell_6t_3 inst_cell_98_118 ( BL118, BLN118, WL98);
sram_cell_6t_3 inst_cell_98_117 ( BL117, BLN117, WL98);
sram_cell_6t_3 inst_cell_98_116 ( BL116, BLN116, WL98);
sram_cell_6t_3 inst_cell_98_115 ( BL115, BLN115, WL98);
sram_cell_6t_3 inst_cell_98_114 ( BL114, BLN114, WL98);
sram_cell_6t_3 inst_cell_98_113 ( BL113, BLN113, WL98);
sram_cell_6t_3 inst_cell_98_112 ( BL112, BLN112, WL98);
sram_cell_6t_3 inst_cell_98_111 ( BL111, BLN111, WL98);
sram_cell_6t_3 inst_cell_98_110 ( BL110, BLN110, WL98);
sram_cell_6t_3 inst_cell_98_109 ( BL109, BLN109, WL98);
sram_cell_6t_3 inst_cell_98_108 ( BL108, BLN108, WL98);
sram_cell_6t_3 inst_cell_98_107 ( BL107, BLN107, WL98);
sram_cell_6t_3 inst_cell_98_106 ( BL106, BLN106, WL98);
sram_cell_6t_3 inst_cell_98_105 ( BL105, BLN105, WL98);
sram_cell_6t_3 inst_cell_98_104 ( BL104, BLN104, WL98);
sram_cell_6t_3 inst_cell_98_103 ( BL103, BLN103, WL98);
sram_cell_6t_3 inst_cell_98_102 ( BL102, BLN102, WL98);
sram_cell_6t_3 inst_cell_98_101 ( BL101, BLN101, WL98);
sram_cell_6t_3 inst_cell_98_100 ( BL100, BLN100, WL98);
sram_cell_6t_3 inst_cell_98_99 ( BL99, BLN99, WL98);
sram_cell_6t_3 inst_cell_98_98 ( BL98, BLN98, WL98);
sram_cell_6t_3 inst_cell_98_97 ( BL97, BLN97, WL98);
sram_cell_6t_3 inst_cell_98_96 ( BL96, BLN96, WL98);
sram_cell_6t_3 inst_cell_98_95 ( BL95, BLN95, WL98);
sram_cell_6t_3 inst_cell_98_94 ( BL94, BLN94, WL98);
sram_cell_6t_3 inst_cell_98_93 ( BL93, BLN93, WL98);
sram_cell_6t_3 inst_cell_98_92 ( BL92, BLN92, WL98);
sram_cell_6t_3 inst_cell_98_91 ( BL91, BLN91, WL98);
sram_cell_6t_3 inst_cell_98_90 ( BL90, BLN90, WL98);
sram_cell_6t_3 inst_cell_98_89 ( BL89, BLN89, WL98);
sram_cell_6t_3 inst_cell_98_88 ( BL88, BLN88, WL98);
sram_cell_6t_3 inst_cell_98_87 ( BL87, BLN87, WL98);
sram_cell_6t_3 inst_cell_98_86 ( BL86, BLN86, WL98);
sram_cell_6t_3 inst_cell_98_85 ( BL85, BLN85, WL98);
sram_cell_6t_3 inst_cell_98_84 ( BL84, BLN84, WL98);
sram_cell_6t_3 inst_cell_98_83 ( BL83, BLN83, WL98);
sram_cell_6t_3 inst_cell_98_82 ( BL82, BLN82, WL98);
sram_cell_6t_3 inst_cell_98_81 ( BL81, BLN81, WL98);
sram_cell_6t_3 inst_cell_98_80 ( BL80, BLN80, WL98);
sram_cell_6t_3 inst_cell_98_79 ( BL79, BLN79, WL98);
sram_cell_6t_3 inst_cell_98_78 ( BL78, BLN78, WL98);
sram_cell_6t_3 inst_cell_98_77 ( BL77, BLN77, WL98);
sram_cell_6t_3 inst_cell_98_76 ( BL76, BLN76, WL98);
sram_cell_6t_3 inst_cell_98_75 ( BL75, BLN75, WL98);
sram_cell_6t_3 inst_cell_98_74 ( BL74, BLN74, WL98);
sram_cell_6t_3 inst_cell_98_73 ( BL73, BLN73, WL98);
sram_cell_6t_3 inst_cell_98_72 ( BL72, BLN72, WL98);
sram_cell_6t_3 inst_cell_98_71 ( BL71, BLN71, WL98);
sram_cell_6t_3 inst_cell_98_70 ( BL70, BLN70, WL98);
sram_cell_6t_3 inst_cell_98_69 ( BL69, BLN69, WL98);
sram_cell_6t_3 inst_cell_98_68 ( BL68, BLN68, WL98);
sram_cell_6t_3 inst_cell_98_67 ( BL67, BLN67, WL98);
sram_cell_6t_3 inst_cell_98_66 ( BL66, BLN66, WL98);
sram_cell_6t_3 inst_cell_98_65 ( BL65, BLN65, WL98);
sram_cell_6t_3 inst_cell_98_64 ( BL64, BLN64, WL98);
sram_cell_6t_3 inst_cell_98_63 ( BL63, BLN63, WL98);
sram_cell_6t_3 inst_cell_98_62 ( BL62, BLN62, WL98);
sram_cell_6t_3 inst_cell_98_61 ( BL61, BLN61, WL98);
sram_cell_6t_3 inst_cell_98_60 ( BL60, BLN60, WL98);
sram_cell_6t_3 inst_cell_98_59 ( BL59, BLN59, WL98);
sram_cell_6t_3 inst_cell_98_58 ( BL58, BLN58, WL98);
sram_cell_6t_3 inst_cell_98_57 ( BL57, BLN57, WL98);
sram_cell_6t_3 inst_cell_98_56 ( BL56, BLN56, WL98);
sram_cell_6t_3 inst_cell_98_55 ( BL55, BLN55, WL98);
sram_cell_6t_3 inst_cell_98_54 ( BL54, BLN54, WL98);
sram_cell_6t_3 inst_cell_98_53 ( BL53, BLN53, WL98);
sram_cell_6t_3 inst_cell_98_52 ( BL52, BLN52, WL98);
sram_cell_6t_3 inst_cell_98_51 ( BL51, BLN51, WL98);
sram_cell_6t_3 inst_cell_98_50 ( BL50, BLN50, WL98);
sram_cell_6t_3 inst_cell_98_49 ( BL49, BLN49, WL98);
sram_cell_6t_3 inst_cell_98_48 ( BL48, BLN48, WL98);
sram_cell_6t_3 inst_cell_98_47 ( BL47, BLN47, WL98);
sram_cell_6t_3 inst_cell_98_46 ( BL46, BLN46, WL98);
sram_cell_6t_3 inst_cell_98_45 ( BL45, BLN45, WL98);
sram_cell_6t_3 inst_cell_98_44 ( BL44, BLN44, WL98);
sram_cell_6t_3 inst_cell_98_43 ( BL43, BLN43, WL98);
sram_cell_6t_3 inst_cell_98_42 ( BL42, BLN42, WL98);
sram_cell_6t_3 inst_cell_98_41 ( BL41, BLN41, WL98);
sram_cell_6t_3 inst_cell_98_40 ( BL40, BLN40, WL98);
sram_cell_6t_3 inst_cell_98_39 ( BL39, BLN39, WL98);
sram_cell_6t_3 inst_cell_98_38 ( BL38, BLN38, WL98);
sram_cell_6t_3 inst_cell_98_37 ( BL37, BLN37, WL98);
sram_cell_6t_3 inst_cell_98_36 ( BL36, BLN36, WL98);
sram_cell_6t_3 inst_cell_98_35 ( BL35, BLN35, WL98);
sram_cell_6t_3 inst_cell_98_34 ( BL34, BLN34, WL98);
sram_cell_6t_3 inst_cell_98_33 ( BL33, BLN33, WL98);
sram_cell_6t_3 inst_cell_98_32 ( BL32, BLN32, WL98);
sram_cell_6t_3 inst_cell_98_31 ( BL31, BLN31, WL98);
sram_cell_6t_3 inst_cell_98_30 ( BL30, BLN30, WL98);
sram_cell_6t_3 inst_cell_98_29 ( BL29, BLN29, WL98);
sram_cell_6t_3 inst_cell_98_28 ( BL28, BLN28, WL98);
sram_cell_6t_3 inst_cell_98_27 ( BL27, BLN27, WL98);
sram_cell_6t_3 inst_cell_98_26 ( BL26, BLN26, WL98);
sram_cell_6t_3 inst_cell_98_25 ( BL25, BLN25, WL98);
sram_cell_6t_3 inst_cell_98_24 ( BL24, BLN24, WL98);
sram_cell_6t_3 inst_cell_98_23 ( BL23, BLN23, WL98);
sram_cell_6t_3 inst_cell_98_22 ( BL22, BLN22, WL98);
sram_cell_6t_3 inst_cell_98_21 ( BL21, BLN21, WL98);
sram_cell_6t_3 inst_cell_98_20 ( BL20, BLN20, WL98);
sram_cell_6t_3 inst_cell_98_19 ( BL19, BLN19, WL98);
sram_cell_6t_3 inst_cell_98_18 ( BL18, BLN18, WL98);
sram_cell_6t_3 inst_cell_98_17 ( BL17, BLN17, WL98);
sram_cell_6t_3 inst_cell_98_16 ( BL16, BLN16, WL98);
sram_cell_6t_3 inst_cell_98_15 ( BL15, BLN15, WL98);
sram_cell_6t_3 inst_cell_98_14 ( BL14, BLN14, WL98);
sram_cell_6t_3 inst_cell_98_13 ( BL13, BLN13, WL98);
sram_cell_6t_3 inst_cell_98_12 ( BL12, BLN12, WL98);
sram_cell_6t_3 inst_cell_98_11 ( BL11, BLN11, WL98);
sram_cell_6t_3 inst_cell_98_10 ( BL10, BLN10, WL98);
sram_cell_6t_3 inst_cell_98_9 ( BL9, BLN9, WL98);
sram_cell_6t_3 inst_cell_98_8 ( BL8, BLN8, WL98);
sram_cell_6t_3 inst_cell_98_7 ( BL7, BLN7, WL98);
sram_cell_6t_3 inst_cell_98_6 ( BL6, BLN6, WL98);
sram_cell_6t_3 inst_cell_98_5 ( BL5, BLN5, WL98);
sram_cell_6t_3 inst_cell_98_4 ( BL4, BLN4, WL98);
sram_cell_6t_3 inst_cell_98_3 ( BL3, BLN3, WL98);
sram_cell_6t_3 inst_cell_98_2 ( BL2, BLN2, WL98);
sram_cell_6t_3 inst_cell_98_1 ( BL1, BLN1, WL98);
sram_cell_6t_3 inst_cell_98_0 ( BL0, BLN0, WL98);
sram_cell_6t_3 inst_cell_97_127 ( BL127, BLN127, WL97);
sram_cell_6t_3 inst_cell_97_126 ( BL126, BLN126, WL97);
sram_cell_6t_3 inst_cell_97_125 ( BL125, BLN125, WL97);
sram_cell_6t_3 inst_cell_97_124 ( BL124, BLN124, WL97);
sram_cell_6t_3 inst_cell_97_123 ( BL123, BLN123, WL97);
sram_cell_6t_3 inst_cell_97_122 ( BL122, BLN122, WL97);
sram_cell_6t_3 inst_cell_97_121 ( BL121, BLN121, WL97);
sram_cell_6t_3 inst_cell_97_120 ( BL120, BLN120, WL97);
sram_cell_6t_3 inst_cell_97_119 ( BL119, BLN119, WL97);
sram_cell_6t_3 inst_cell_97_118 ( BL118, BLN118, WL97);
sram_cell_6t_3 inst_cell_97_117 ( BL117, BLN117, WL97);
sram_cell_6t_3 inst_cell_97_116 ( BL116, BLN116, WL97);
sram_cell_6t_3 inst_cell_97_115 ( BL115, BLN115, WL97);
sram_cell_6t_3 inst_cell_97_114 ( BL114, BLN114, WL97);
sram_cell_6t_3 inst_cell_97_113 ( BL113, BLN113, WL97);
sram_cell_6t_3 inst_cell_97_112 ( BL112, BLN112, WL97);
sram_cell_6t_3 inst_cell_97_111 ( BL111, BLN111, WL97);
sram_cell_6t_3 inst_cell_97_110 ( BL110, BLN110, WL97);
sram_cell_6t_3 inst_cell_97_109 ( BL109, BLN109, WL97);
sram_cell_6t_3 inst_cell_97_108 ( BL108, BLN108, WL97);
sram_cell_6t_3 inst_cell_97_107 ( BL107, BLN107, WL97);
sram_cell_6t_3 inst_cell_97_106 ( BL106, BLN106, WL97);
sram_cell_6t_3 inst_cell_97_105 ( BL105, BLN105, WL97);
sram_cell_6t_3 inst_cell_97_104 ( BL104, BLN104, WL97);
sram_cell_6t_3 inst_cell_97_103 ( BL103, BLN103, WL97);
sram_cell_6t_3 inst_cell_97_102 ( BL102, BLN102, WL97);
sram_cell_6t_3 inst_cell_97_101 ( BL101, BLN101, WL97);
sram_cell_6t_3 inst_cell_97_100 ( BL100, BLN100, WL97);
sram_cell_6t_3 inst_cell_97_99 ( BL99, BLN99, WL97);
sram_cell_6t_3 inst_cell_97_98 ( BL98, BLN98, WL97);
sram_cell_6t_3 inst_cell_97_97 ( BL97, BLN97, WL97);
sram_cell_6t_3 inst_cell_97_96 ( BL96, BLN96, WL97);
sram_cell_6t_3 inst_cell_97_95 ( BL95, BLN95, WL97);
sram_cell_6t_3 inst_cell_97_94 ( BL94, BLN94, WL97);
sram_cell_6t_3 inst_cell_97_93 ( BL93, BLN93, WL97);
sram_cell_6t_3 inst_cell_97_92 ( BL92, BLN92, WL97);
sram_cell_6t_3 inst_cell_97_91 ( BL91, BLN91, WL97);
sram_cell_6t_3 inst_cell_97_90 ( BL90, BLN90, WL97);
sram_cell_6t_3 inst_cell_97_89 ( BL89, BLN89, WL97);
sram_cell_6t_3 inst_cell_97_88 ( BL88, BLN88, WL97);
sram_cell_6t_3 inst_cell_97_87 ( BL87, BLN87, WL97);
sram_cell_6t_3 inst_cell_97_86 ( BL86, BLN86, WL97);
sram_cell_6t_3 inst_cell_97_85 ( BL85, BLN85, WL97);
sram_cell_6t_3 inst_cell_97_84 ( BL84, BLN84, WL97);
sram_cell_6t_3 inst_cell_97_83 ( BL83, BLN83, WL97);
sram_cell_6t_3 inst_cell_97_82 ( BL82, BLN82, WL97);
sram_cell_6t_3 inst_cell_97_81 ( BL81, BLN81, WL97);
sram_cell_6t_3 inst_cell_97_80 ( BL80, BLN80, WL97);
sram_cell_6t_3 inst_cell_97_79 ( BL79, BLN79, WL97);
sram_cell_6t_3 inst_cell_97_78 ( BL78, BLN78, WL97);
sram_cell_6t_3 inst_cell_97_77 ( BL77, BLN77, WL97);
sram_cell_6t_3 inst_cell_97_76 ( BL76, BLN76, WL97);
sram_cell_6t_3 inst_cell_97_75 ( BL75, BLN75, WL97);
sram_cell_6t_3 inst_cell_97_74 ( BL74, BLN74, WL97);
sram_cell_6t_3 inst_cell_97_73 ( BL73, BLN73, WL97);
sram_cell_6t_3 inst_cell_97_72 ( BL72, BLN72, WL97);
sram_cell_6t_3 inst_cell_97_71 ( BL71, BLN71, WL97);
sram_cell_6t_3 inst_cell_97_70 ( BL70, BLN70, WL97);
sram_cell_6t_3 inst_cell_97_69 ( BL69, BLN69, WL97);
sram_cell_6t_3 inst_cell_97_68 ( BL68, BLN68, WL97);
sram_cell_6t_3 inst_cell_97_67 ( BL67, BLN67, WL97);
sram_cell_6t_3 inst_cell_97_66 ( BL66, BLN66, WL97);
sram_cell_6t_3 inst_cell_97_65 ( BL65, BLN65, WL97);
sram_cell_6t_3 inst_cell_97_64 ( BL64, BLN64, WL97);
sram_cell_6t_3 inst_cell_97_63 ( BL63, BLN63, WL97);
sram_cell_6t_3 inst_cell_97_62 ( BL62, BLN62, WL97);
sram_cell_6t_3 inst_cell_97_61 ( BL61, BLN61, WL97);
sram_cell_6t_3 inst_cell_97_60 ( BL60, BLN60, WL97);
sram_cell_6t_3 inst_cell_97_59 ( BL59, BLN59, WL97);
sram_cell_6t_3 inst_cell_97_58 ( BL58, BLN58, WL97);
sram_cell_6t_3 inst_cell_97_57 ( BL57, BLN57, WL97);
sram_cell_6t_3 inst_cell_97_56 ( BL56, BLN56, WL97);
sram_cell_6t_3 inst_cell_97_55 ( BL55, BLN55, WL97);
sram_cell_6t_3 inst_cell_97_54 ( BL54, BLN54, WL97);
sram_cell_6t_3 inst_cell_97_53 ( BL53, BLN53, WL97);
sram_cell_6t_3 inst_cell_97_52 ( BL52, BLN52, WL97);
sram_cell_6t_3 inst_cell_97_51 ( BL51, BLN51, WL97);
sram_cell_6t_3 inst_cell_97_50 ( BL50, BLN50, WL97);
sram_cell_6t_3 inst_cell_97_49 ( BL49, BLN49, WL97);
sram_cell_6t_3 inst_cell_97_48 ( BL48, BLN48, WL97);
sram_cell_6t_3 inst_cell_97_47 ( BL47, BLN47, WL97);
sram_cell_6t_3 inst_cell_97_46 ( BL46, BLN46, WL97);
sram_cell_6t_3 inst_cell_97_45 ( BL45, BLN45, WL97);
sram_cell_6t_3 inst_cell_97_44 ( BL44, BLN44, WL97);
sram_cell_6t_3 inst_cell_97_43 ( BL43, BLN43, WL97);
sram_cell_6t_3 inst_cell_97_42 ( BL42, BLN42, WL97);
sram_cell_6t_3 inst_cell_97_41 ( BL41, BLN41, WL97);
sram_cell_6t_3 inst_cell_97_40 ( BL40, BLN40, WL97);
sram_cell_6t_3 inst_cell_97_39 ( BL39, BLN39, WL97);
sram_cell_6t_3 inst_cell_97_38 ( BL38, BLN38, WL97);
sram_cell_6t_3 inst_cell_97_37 ( BL37, BLN37, WL97);
sram_cell_6t_3 inst_cell_97_36 ( BL36, BLN36, WL97);
sram_cell_6t_3 inst_cell_97_35 ( BL35, BLN35, WL97);
sram_cell_6t_3 inst_cell_97_34 ( BL34, BLN34, WL97);
sram_cell_6t_3 inst_cell_97_33 ( BL33, BLN33, WL97);
sram_cell_6t_3 inst_cell_97_32 ( BL32, BLN32, WL97);
sram_cell_6t_3 inst_cell_97_31 ( BL31, BLN31, WL97);
sram_cell_6t_3 inst_cell_97_30 ( BL30, BLN30, WL97);
sram_cell_6t_3 inst_cell_97_29 ( BL29, BLN29, WL97);
sram_cell_6t_3 inst_cell_97_28 ( BL28, BLN28, WL97);
sram_cell_6t_3 inst_cell_97_27 ( BL27, BLN27, WL97);
sram_cell_6t_3 inst_cell_97_26 ( BL26, BLN26, WL97);
sram_cell_6t_3 inst_cell_97_25 ( BL25, BLN25, WL97);
sram_cell_6t_3 inst_cell_97_24 ( BL24, BLN24, WL97);
sram_cell_6t_3 inst_cell_97_23 ( BL23, BLN23, WL97);
sram_cell_6t_3 inst_cell_97_22 ( BL22, BLN22, WL97);
sram_cell_6t_3 inst_cell_97_21 ( BL21, BLN21, WL97);
sram_cell_6t_3 inst_cell_97_20 ( BL20, BLN20, WL97);
sram_cell_6t_3 inst_cell_97_19 ( BL19, BLN19, WL97);
sram_cell_6t_3 inst_cell_97_18 ( BL18, BLN18, WL97);
sram_cell_6t_3 inst_cell_97_17 ( BL17, BLN17, WL97);
sram_cell_6t_3 inst_cell_97_16 ( BL16, BLN16, WL97);
sram_cell_6t_3 inst_cell_97_15 ( BL15, BLN15, WL97);
sram_cell_6t_3 inst_cell_97_14 ( BL14, BLN14, WL97);
sram_cell_6t_3 inst_cell_97_13 ( BL13, BLN13, WL97);
sram_cell_6t_3 inst_cell_97_12 ( BL12, BLN12, WL97);
sram_cell_6t_3 inst_cell_97_11 ( BL11, BLN11, WL97);
sram_cell_6t_3 inst_cell_97_10 ( BL10, BLN10, WL97);
sram_cell_6t_3 inst_cell_97_9 ( BL9, BLN9, WL97);
sram_cell_6t_3 inst_cell_97_8 ( BL8, BLN8, WL97);
sram_cell_6t_3 inst_cell_97_7 ( BL7, BLN7, WL97);
sram_cell_6t_3 inst_cell_97_6 ( BL6, BLN6, WL97);
sram_cell_6t_3 inst_cell_97_5 ( BL5, BLN5, WL97);
sram_cell_6t_3 inst_cell_97_4 ( BL4, BLN4, WL97);
sram_cell_6t_3 inst_cell_97_3 ( BL3, BLN3, WL97);
sram_cell_6t_3 inst_cell_97_2 ( BL2, BLN2, WL97);
sram_cell_6t_3 inst_cell_97_1 ( BL1, BLN1, WL97);
sram_cell_6t_3 inst_cell_97_0 ( BL0, BLN0, WL97);
sram_cell_6t_3 inst_cell_96_127 ( BL127, BLN127, WL96);
sram_cell_6t_3 inst_cell_96_126 ( BL126, BLN126, WL96);
sram_cell_6t_3 inst_cell_96_125 ( BL125, BLN125, WL96);
sram_cell_6t_3 inst_cell_96_124 ( BL124, BLN124, WL96);
sram_cell_6t_3 inst_cell_96_123 ( BL123, BLN123, WL96);
sram_cell_6t_3 inst_cell_96_122 ( BL122, BLN122, WL96);
sram_cell_6t_3 inst_cell_96_121 ( BL121, BLN121, WL96);
sram_cell_6t_3 inst_cell_96_120 ( BL120, BLN120, WL96);
sram_cell_6t_3 inst_cell_96_119 ( BL119, BLN119, WL96);
sram_cell_6t_3 inst_cell_96_118 ( BL118, BLN118, WL96);
sram_cell_6t_3 inst_cell_96_117 ( BL117, BLN117, WL96);
sram_cell_6t_3 inst_cell_96_116 ( BL116, BLN116, WL96);
sram_cell_6t_3 inst_cell_96_115 ( BL115, BLN115, WL96);
sram_cell_6t_3 inst_cell_96_114 ( BL114, BLN114, WL96);
sram_cell_6t_3 inst_cell_96_113 ( BL113, BLN113, WL96);
sram_cell_6t_3 inst_cell_96_112 ( BL112, BLN112, WL96);
sram_cell_6t_3 inst_cell_96_111 ( BL111, BLN111, WL96);
sram_cell_6t_3 inst_cell_96_110 ( BL110, BLN110, WL96);
sram_cell_6t_3 inst_cell_96_109 ( BL109, BLN109, WL96);
sram_cell_6t_3 inst_cell_96_108 ( BL108, BLN108, WL96);
sram_cell_6t_3 inst_cell_96_107 ( BL107, BLN107, WL96);
sram_cell_6t_3 inst_cell_96_106 ( BL106, BLN106, WL96);
sram_cell_6t_3 inst_cell_96_105 ( BL105, BLN105, WL96);
sram_cell_6t_3 inst_cell_96_104 ( BL104, BLN104, WL96);
sram_cell_6t_3 inst_cell_96_103 ( BL103, BLN103, WL96);
sram_cell_6t_3 inst_cell_96_102 ( BL102, BLN102, WL96);
sram_cell_6t_3 inst_cell_96_101 ( BL101, BLN101, WL96);
sram_cell_6t_3 inst_cell_96_100 ( BL100, BLN100, WL96);
sram_cell_6t_3 inst_cell_96_99 ( BL99, BLN99, WL96);
sram_cell_6t_3 inst_cell_96_98 ( BL98, BLN98, WL96);
sram_cell_6t_3 inst_cell_96_97 ( BL97, BLN97, WL96);
sram_cell_6t_3 inst_cell_96_96 ( BL96, BLN96, WL96);
sram_cell_6t_3 inst_cell_96_95 ( BL95, BLN95, WL96);
sram_cell_6t_3 inst_cell_96_94 ( BL94, BLN94, WL96);
sram_cell_6t_3 inst_cell_96_93 ( BL93, BLN93, WL96);
sram_cell_6t_3 inst_cell_96_92 ( BL92, BLN92, WL96);
sram_cell_6t_3 inst_cell_96_91 ( BL91, BLN91, WL96);
sram_cell_6t_3 inst_cell_96_90 ( BL90, BLN90, WL96);
sram_cell_6t_3 inst_cell_96_89 ( BL89, BLN89, WL96);
sram_cell_6t_3 inst_cell_96_88 ( BL88, BLN88, WL96);
sram_cell_6t_3 inst_cell_96_87 ( BL87, BLN87, WL96);
sram_cell_6t_3 inst_cell_96_86 ( BL86, BLN86, WL96);
sram_cell_6t_3 inst_cell_96_85 ( BL85, BLN85, WL96);
sram_cell_6t_3 inst_cell_96_84 ( BL84, BLN84, WL96);
sram_cell_6t_3 inst_cell_96_83 ( BL83, BLN83, WL96);
sram_cell_6t_3 inst_cell_96_82 ( BL82, BLN82, WL96);
sram_cell_6t_3 inst_cell_96_81 ( BL81, BLN81, WL96);
sram_cell_6t_3 inst_cell_96_80 ( BL80, BLN80, WL96);
sram_cell_6t_3 inst_cell_96_79 ( BL79, BLN79, WL96);
sram_cell_6t_3 inst_cell_96_78 ( BL78, BLN78, WL96);
sram_cell_6t_3 inst_cell_96_77 ( BL77, BLN77, WL96);
sram_cell_6t_3 inst_cell_96_76 ( BL76, BLN76, WL96);
sram_cell_6t_3 inst_cell_96_75 ( BL75, BLN75, WL96);
sram_cell_6t_3 inst_cell_96_74 ( BL74, BLN74, WL96);
sram_cell_6t_3 inst_cell_96_73 ( BL73, BLN73, WL96);
sram_cell_6t_3 inst_cell_96_72 ( BL72, BLN72, WL96);
sram_cell_6t_3 inst_cell_96_71 ( BL71, BLN71, WL96);
sram_cell_6t_3 inst_cell_96_70 ( BL70, BLN70, WL96);
sram_cell_6t_3 inst_cell_96_69 ( BL69, BLN69, WL96);
sram_cell_6t_3 inst_cell_96_68 ( BL68, BLN68, WL96);
sram_cell_6t_3 inst_cell_96_67 ( BL67, BLN67, WL96);
sram_cell_6t_3 inst_cell_96_66 ( BL66, BLN66, WL96);
sram_cell_6t_3 inst_cell_96_65 ( BL65, BLN65, WL96);
sram_cell_6t_3 inst_cell_96_64 ( BL64, BLN64, WL96);
sram_cell_6t_3 inst_cell_96_63 ( BL63, BLN63, WL96);
sram_cell_6t_3 inst_cell_96_62 ( BL62, BLN62, WL96);
sram_cell_6t_3 inst_cell_96_61 ( BL61, BLN61, WL96);
sram_cell_6t_3 inst_cell_96_60 ( BL60, BLN60, WL96);
sram_cell_6t_3 inst_cell_96_59 ( BL59, BLN59, WL96);
sram_cell_6t_3 inst_cell_96_58 ( BL58, BLN58, WL96);
sram_cell_6t_3 inst_cell_96_57 ( BL57, BLN57, WL96);
sram_cell_6t_3 inst_cell_96_56 ( BL56, BLN56, WL96);
sram_cell_6t_3 inst_cell_96_55 ( BL55, BLN55, WL96);
sram_cell_6t_3 inst_cell_96_54 ( BL54, BLN54, WL96);
sram_cell_6t_3 inst_cell_96_53 ( BL53, BLN53, WL96);
sram_cell_6t_3 inst_cell_96_52 ( BL52, BLN52, WL96);
sram_cell_6t_3 inst_cell_96_51 ( BL51, BLN51, WL96);
sram_cell_6t_3 inst_cell_96_50 ( BL50, BLN50, WL96);
sram_cell_6t_3 inst_cell_96_49 ( BL49, BLN49, WL96);
sram_cell_6t_3 inst_cell_96_48 ( BL48, BLN48, WL96);
sram_cell_6t_3 inst_cell_96_47 ( BL47, BLN47, WL96);
sram_cell_6t_3 inst_cell_96_46 ( BL46, BLN46, WL96);
sram_cell_6t_3 inst_cell_96_45 ( BL45, BLN45, WL96);
sram_cell_6t_3 inst_cell_96_44 ( BL44, BLN44, WL96);
sram_cell_6t_3 inst_cell_96_43 ( BL43, BLN43, WL96);
sram_cell_6t_3 inst_cell_96_42 ( BL42, BLN42, WL96);
sram_cell_6t_3 inst_cell_96_41 ( BL41, BLN41, WL96);
sram_cell_6t_3 inst_cell_96_40 ( BL40, BLN40, WL96);
sram_cell_6t_3 inst_cell_96_39 ( BL39, BLN39, WL96);
sram_cell_6t_3 inst_cell_96_38 ( BL38, BLN38, WL96);
sram_cell_6t_3 inst_cell_96_37 ( BL37, BLN37, WL96);
sram_cell_6t_3 inst_cell_96_36 ( BL36, BLN36, WL96);
sram_cell_6t_3 inst_cell_96_35 ( BL35, BLN35, WL96);
sram_cell_6t_3 inst_cell_96_34 ( BL34, BLN34, WL96);
sram_cell_6t_3 inst_cell_96_33 ( BL33, BLN33, WL96);
sram_cell_6t_3 inst_cell_96_32 ( BL32, BLN32, WL96);
sram_cell_6t_3 inst_cell_96_31 ( BL31, BLN31, WL96);
sram_cell_6t_3 inst_cell_96_30 ( BL30, BLN30, WL96);
sram_cell_6t_3 inst_cell_96_29 ( BL29, BLN29, WL96);
sram_cell_6t_3 inst_cell_96_28 ( BL28, BLN28, WL96);
sram_cell_6t_3 inst_cell_96_27 ( BL27, BLN27, WL96);
sram_cell_6t_3 inst_cell_96_26 ( BL26, BLN26, WL96);
sram_cell_6t_3 inst_cell_96_25 ( BL25, BLN25, WL96);
sram_cell_6t_3 inst_cell_96_24 ( BL24, BLN24, WL96);
sram_cell_6t_3 inst_cell_96_23 ( BL23, BLN23, WL96);
sram_cell_6t_3 inst_cell_96_22 ( BL22, BLN22, WL96);
sram_cell_6t_3 inst_cell_96_21 ( BL21, BLN21, WL96);
sram_cell_6t_3 inst_cell_96_20 ( BL20, BLN20, WL96);
sram_cell_6t_3 inst_cell_96_19 ( BL19, BLN19, WL96);
sram_cell_6t_3 inst_cell_96_18 ( BL18, BLN18, WL96);
sram_cell_6t_3 inst_cell_96_17 ( BL17, BLN17, WL96);
sram_cell_6t_3 inst_cell_96_16 ( BL16, BLN16, WL96);
sram_cell_6t_3 inst_cell_96_15 ( BL15, BLN15, WL96);
sram_cell_6t_3 inst_cell_96_14 ( BL14, BLN14, WL96);
sram_cell_6t_3 inst_cell_96_13 ( BL13, BLN13, WL96);
sram_cell_6t_3 inst_cell_96_12 ( BL12, BLN12, WL96);
sram_cell_6t_3 inst_cell_96_11 ( BL11, BLN11, WL96);
sram_cell_6t_3 inst_cell_96_10 ( BL10, BLN10, WL96);
sram_cell_6t_3 inst_cell_96_9 ( BL9, BLN9, WL96);
sram_cell_6t_3 inst_cell_96_8 ( BL8, BLN8, WL96);
sram_cell_6t_3 inst_cell_96_7 ( BL7, BLN7, WL96);
sram_cell_6t_3 inst_cell_96_6 ( BL6, BLN6, WL96);
sram_cell_6t_3 inst_cell_96_5 ( BL5, BLN5, WL96);
sram_cell_6t_3 inst_cell_96_4 ( BL4, BLN4, WL96);
sram_cell_6t_3 inst_cell_96_3 ( BL3, BLN3, WL96);
sram_cell_6t_3 inst_cell_96_2 ( BL2, BLN2, WL96);
sram_cell_6t_3 inst_cell_96_1 ( BL1, BLN1, WL96);
sram_cell_6t_3 inst_cell_96_0 ( BL0, BLN0, WL96);
sram_cell_6t_3 inst_cell_95_127 ( BL127, BLN127, WL95);
sram_cell_6t_3 inst_cell_95_126 ( BL126, BLN126, WL95);
sram_cell_6t_3 inst_cell_95_125 ( BL125, BLN125, WL95);
sram_cell_6t_3 inst_cell_95_124 ( BL124, BLN124, WL95);
sram_cell_6t_3 inst_cell_95_123 ( BL123, BLN123, WL95);
sram_cell_6t_3 inst_cell_95_122 ( BL122, BLN122, WL95);
sram_cell_6t_3 inst_cell_95_121 ( BL121, BLN121, WL95);
sram_cell_6t_3 inst_cell_95_120 ( BL120, BLN120, WL95);
sram_cell_6t_3 inst_cell_95_119 ( BL119, BLN119, WL95);
sram_cell_6t_3 inst_cell_95_118 ( BL118, BLN118, WL95);
sram_cell_6t_3 inst_cell_95_117 ( BL117, BLN117, WL95);
sram_cell_6t_3 inst_cell_95_116 ( BL116, BLN116, WL95);
sram_cell_6t_3 inst_cell_95_115 ( BL115, BLN115, WL95);
sram_cell_6t_3 inst_cell_95_114 ( BL114, BLN114, WL95);
sram_cell_6t_3 inst_cell_95_113 ( BL113, BLN113, WL95);
sram_cell_6t_3 inst_cell_95_112 ( BL112, BLN112, WL95);
sram_cell_6t_3 inst_cell_95_111 ( BL111, BLN111, WL95);
sram_cell_6t_3 inst_cell_95_110 ( BL110, BLN110, WL95);
sram_cell_6t_3 inst_cell_95_109 ( BL109, BLN109, WL95);
sram_cell_6t_3 inst_cell_95_108 ( BL108, BLN108, WL95);
sram_cell_6t_3 inst_cell_95_107 ( BL107, BLN107, WL95);
sram_cell_6t_3 inst_cell_95_106 ( BL106, BLN106, WL95);
sram_cell_6t_3 inst_cell_95_105 ( BL105, BLN105, WL95);
sram_cell_6t_3 inst_cell_95_104 ( BL104, BLN104, WL95);
sram_cell_6t_3 inst_cell_95_103 ( BL103, BLN103, WL95);
sram_cell_6t_3 inst_cell_95_102 ( BL102, BLN102, WL95);
sram_cell_6t_3 inst_cell_95_101 ( BL101, BLN101, WL95);
sram_cell_6t_3 inst_cell_95_100 ( BL100, BLN100, WL95);
sram_cell_6t_3 inst_cell_95_99 ( BL99, BLN99, WL95);
sram_cell_6t_3 inst_cell_95_98 ( BL98, BLN98, WL95);
sram_cell_6t_3 inst_cell_95_97 ( BL97, BLN97, WL95);
sram_cell_6t_3 inst_cell_95_96 ( BL96, BLN96, WL95);
sram_cell_6t_3 inst_cell_95_95 ( BL95, BLN95, WL95);
sram_cell_6t_3 inst_cell_95_94 ( BL94, BLN94, WL95);
sram_cell_6t_3 inst_cell_95_93 ( BL93, BLN93, WL95);
sram_cell_6t_3 inst_cell_95_92 ( BL92, BLN92, WL95);
sram_cell_6t_3 inst_cell_95_91 ( BL91, BLN91, WL95);
sram_cell_6t_3 inst_cell_95_90 ( BL90, BLN90, WL95);
sram_cell_6t_3 inst_cell_95_89 ( BL89, BLN89, WL95);
sram_cell_6t_3 inst_cell_95_88 ( BL88, BLN88, WL95);
sram_cell_6t_3 inst_cell_95_87 ( BL87, BLN87, WL95);
sram_cell_6t_3 inst_cell_95_86 ( BL86, BLN86, WL95);
sram_cell_6t_3 inst_cell_95_85 ( BL85, BLN85, WL95);
sram_cell_6t_3 inst_cell_95_84 ( BL84, BLN84, WL95);
sram_cell_6t_3 inst_cell_95_83 ( BL83, BLN83, WL95);
sram_cell_6t_3 inst_cell_95_82 ( BL82, BLN82, WL95);
sram_cell_6t_3 inst_cell_95_81 ( BL81, BLN81, WL95);
sram_cell_6t_3 inst_cell_95_80 ( BL80, BLN80, WL95);
sram_cell_6t_3 inst_cell_95_79 ( BL79, BLN79, WL95);
sram_cell_6t_3 inst_cell_95_78 ( BL78, BLN78, WL95);
sram_cell_6t_3 inst_cell_95_77 ( BL77, BLN77, WL95);
sram_cell_6t_3 inst_cell_95_76 ( BL76, BLN76, WL95);
sram_cell_6t_3 inst_cell_95_75 ( BL75, BLN75, WL95);
sram_cell_6t_3 inst_cell_95_74 ( BL74, BLN74, WL95);
sram_cell_6t_3 inst_cell_95_73 ( BL73, BLN73, WL95);
sram_cell_6t_3 inst_cell_95_72 ( BL72, BLN72, WL95);
sram_cell_6t_3 inst_cell_95_71 ( BL71, BLN71, WL95);
sram_cell_6t_3 inst_cell_95_70 ( BL70, BLN70, WL95);
sram_cell_6t_3 inst_cell_95_69 ( BL69, BLN69, WL95);
sram_cell_6t_3 inst_cell_95_68 ( BL68, BLN68, WL95);
sram_cell_6t_3 inst_cell_95_67 ( BL67, BLN67, WL95);
sram_cell_6t_3 inst_cell_95_66 ( BL66, BLN66, WL95);
sram_cell_6t_3 inst_cell_95_65 ( BL65, BLN65, WL95);
sram_cell_6t_3 inst_cell_95_64 ( BL64, BLN64, WL95);
sram_cell_6t_3 inst_cell_95_63 ( BL63, BLN63, WL95);
sram_cell_6t_3 inst_cell_95_62 ( BL62, BLN62, WL95);
sram_cell_6t_3 inst_cell_95_61 ( BL61, BLN61, WL95);
sram_cell_6t_3 inst_cell_95_60 ( BL60, BLN60, WL95);
sram_cell_6t_3 inst_cell_95_59 ( BL59, BLN59, WL95);
sram_cell_6t_3 inst_cell_95_58 ( BL58, BLN58, WL95);
sram_cell_6t_3 inst_cell_95_57 ( BL57, BLN57, WL95);
sram_cell_6t_3 inst_cell_95_56 ( BL56, BLN56, WL95);
sram_cell_6t_3 inst_cell_95_55 ( BL55, BLN55, WL95);
sram_cell_6t_3 inst_cell_95_54 ( BL54, BLN54, WL95);
sram_cell_6t_3 inst_cell_95_53 ( BL53, BLN53, WL95);
sram_cell_6t_3 inst_cell_95_52 ( BL52, BLN52, WL95);
sram_cell_6t_3 inst_cell_95_51 ( BL51, BLN51, WL95);
sram_cell_6t_3 inst_cell_95_50 ( BL50, BLN50, WL95);
sram_cell_6t_3 inst_cell_95_49 ( BL49, BLN49, WL95);
sram_cell_6t_3 inst_cell_95_48 ( BL48, BLN48, WL95);
sram_cell_6t_3 inst_cell_95_47 ( BL47, BLN47, WL95);
sram_cell_6t_3 inst_cell_95_46 ( BL46, BLN46, WL95);
sram_cell_6t_3 inst_cell_95_45 ( BL45, BLN45, WL95);
sram_cell_6t_3 inst_cell_95_44 ( BL44, BLN44, WL95);
sram_cell_6t_3 inst_cell_95_43 ( BL43, BLN43, WL95);
sram_cell_6t_3 inst_cell_95_42 ( BL42, BLN42, WL95);
sram_cell_6t_3 inst_cell_95_41 ( BL41, BLN41, WL95);
sram_cell_6t_3 inst_cell_95_40 ( BL40, BLN40, WL95);
sram_cell_6t_3 inst_cell_95_39 ( BL39, BLN39, WL95);
sram_cell_6t_3 inst_cell_95_38 ( BL38, BLN38, WL95);
sram_cell_6t_3 inst_cell_95_37 ( BL37, BLN37, WL95);
sram_cell_6t_3 inst_cell_95_36 ( BL36, BLN36, WL95);
sram_cell_6t_3 inst_cell_95_35 ( BL35, BLN35, WL95);
sram_cell_6t_3 inst_cell_95_34 ( BL34, BLN34, WL95);
sram_cell_6t_3 inst_cell_95_33 ( BL33, BLN33, WL95);
sram_cell_6t_3 inst_cell_95_32 ( BL32, BLN32, WL95);
sram_cell_6t_3 inst_cell_95_31 ( BL31, BLN31, WL95);
sram_cell_6t_3 inst_cell_95_30 ( BL30, BLN30, WL95);
sram_cell_6t_3 inst_cell_95_29 ( BL29, BLN29, WL95);
sram_cell_6t_3 inst_cell_95_28 ( BL28, BLN28, WL95);
sram_cell_6t_3 inst_cell_95_27 ( BL27, BLN27, WL95);
sram_cell_6t_3 inst_cell_95_26 ( BL26, BLN26, WL95);
sram_cell_6t_3 inst_cell_95_25 ( BL25, BLN25, WL95);
sram_cell_6t_3 inst_cell_95_24 ( BL24, BLN24, WL95);
sram_cell_6t_3 inst_cell_95_23 ( BL23, BLN23, WL95);
sram_cell_6t_3 inst_cell_95_22 ( BL22, BLN22, WL95);
sram_cell_6t_3 inst_cell_95_21 ( BL21, BLN21, WL95);
sram_cell_6t_3 inst_cell_95_20 ( BL20, BLN20, WL95);
sram_cell_6t_3 inst_cell_95_19 ( BL19, BLN19, WL95);
sram_cell_6t_3 inst_cell_95_18 ( BL18, BLN18, WL95);
sram_cell_6t_3 inst_cell_95_17 ( BL17, BLN17, WL95);
sram_cell_6t_3 inst_cell_95_16 ( BL16, BLN16, WL95);
sram_cell_6t_3 inst_cell_95_15 ( BL15, BLN15, WL95);
sram_cell_6t_3 inst_cell_95_14 ( BL14, BLN14, WL95);
sram_cell_6t_3 inst_cell_95_13 ( BL13, BLN13, WL95);
sram_cell_6t_3 inst_cell_95_12 ( BL12, BLN12, WL95);
sram_cell_6t_3 inst_cell_95_11 ( BL11, BLN11, WL95);
sram_cell_6t_3 inst_cell_95_10 ( BL10, BLN10, WL95);
sram_cell_6t_3 inst_cell_95_9 ( BL9, BLN9, WL95);
sram_cell_6t_3 inst_cell_95_8 ( BL8, BLN8, WL95);
sram_cell_6t_3 inst_cell_95_7 ( BL7, BLN7, WL95);
sram_cell_6t_3 inst_cell_95_6 ( BL6, BLN6, WL95);
sram_cell_6t_3 inst_cell_95_5 ( BL5, BLN5, WL95);
sram_cell_6t_3 inst_cell_95_4 ( BL4, BLN4, WL95);
sram_cell_6t_3 inst_cell_95_3 ( BL3, BLN3, WL95);
sram_cell_6t_3 inst_cell_95_2 ( BL2, BLN2, WL95);
sram_cell_6t_3 inst_cell_95_1 ( BL1, BLN1, WL95);
sram_cell_6t_3 inst_cell_95_0 ( BL0, BLN0, WL95);
sram_cell_6t_3 inst_cell_94_127 ( BL127, BLN127, WL94);
sram_cell_6t_3 inst_cell_94_126 ( BL126, BLN126, WL94);
sram_cell_6t_3 inst_cell_94_125 ( BL125, BLN125, WL94);
sram_cell_6t_3 inst_cell_94_124 ( BL124, BLN124, WL94);
sram_cell_6t_3 inst_cell_94_123 ( BL123, BLN123, WL94);
sram_cell_6t_3 inst_cell_94_122 ( BL122, BLN122, WL94);
sram_cell_6t_3 inst_cell_94_121 ( BL121, BLN121, WL94);
sram_cell_6t_3 inst_cell_94_120 ( BL120, BLN120, WL94);
sram_cell_6t_3 inst_cell_94_119 ( BL119, BLN119, WL94);
sram_cell_6t_3 inst_cell_94_118 ( BL118, BLN118, WL94);
sram_cell_6t_3 inst_cell_94_117 ( BL117, BLN117, WL94);
sram_cell_6t_3 inst_cell_94_116 ( BL116, BLN116, WL94);
sram_cell_6t_3 inst_cell_94_115 ( BL115, BLN115, WL94);
sram_cell_6t_3 inst_cell_94_114 ( BL114, BLN114, WL94);
sram_cell_6t_3 inst_cell_94_113 ( BL113, BLN113, WL94);
sram_cell_6t_3 inst_cell_94_112 ( BL112, BLN112, WL94);
sram_cell_6t_3 inst_cell_94_111 ( BL111, BLN111, WL94);
sram_cell_6t_3 inst_cell_94_110 ( BL110, BLN110, WL94);
sram_cell_6t_3 inst_cell_94_109 ( BL109, BLN109, WL94);
sram_cell_6t_3 inst_cell_94_108 ( BL108, BLN108, WL94);
sram_cell_6t_3 inst_cell_94_107 ( BL107, BLN107, WL94);
sram_cell_6t_3 inst_cell_94_106 ( BL106, BLN106, WL94);
sram_cell_6t_3 inst_cell_94_105 ( BL105, BLN105, WL94);
sram_cell_6t_3 inst_cell_94_104 ( BL104, BLN104, WL94);
sram_cell_6t_3 inst_cell_94_103 ( BL103, BLN103, WL94);
sram_cell_6t_3 inst_cell_94_102 ( BL102, BLN102, WL94);
sram_cell_6t_3 inst_cell_94_101 ( BL101, BLN101, WL94);
sram_cell_6t_3 inst_cell_94_100 ( BL100, BLN100, WL94);
sram_cell_6t_3 inst_cell_94_99 ( BL99, BLN99, WL94);
sram_cell_6t_3 inst_cell_94_98 ( BL98, BLN98, WL94);
sram_cell_6t_3 inst_cell_94_97 ( BL97, BLN97, WL94);
sram_cell_6t_3 inst_cell_94_96 ( BL96, BLN96, WL94);
sram_cell_6t_3 inst_cell_94_95 ( BL95, BLN95, WL94);
sram_cell_6t_3 inst_cell_94_94 ( BL94, BLN94, WL94);
sram_cell_6t_3 inst_cell_94_93 ( BL93, BLN93, WL94);
sram_cell_6t_3 inst_cell_94_92 ( BL92, BLN92, WL94);
sram_cell_6t_3 inst_cell_94_91 ( BL91, BLN91, WL94);
sram_cell_6t_3 inst_cell_94_90 ( BL90, BLN90, WL94);
sram_cell_6t_3 inst_cell_94_89 ( BL89, BLN89, WL94);
sram_cell_6t_3 inst_cell_94_88 ( BL88, BLN88, WL94);
sram_cell_6t_3 inst_cell_94_87 ( BL87, BLN87, WL94);
sram_cell_6t_3 inst_cell_94_86 ( BL86, BLN86, WL94);
sram_cell_6t_3 inst_cell_94_85 ( BL85, BLN85, WL94);
sram_cell_6t_3 inst_cell_94_84 ( BL84, BLN84, WL94);
sram_cell_6t_3 inst_cell_94_83 ( BL83, BLN83, WL94);
sram_cell_6t_3 inst_cell_94_82 ( BL82, BLN82, WL94);
sram_cell_6t_3 inst_cell_94_81 ( BL81, BLN81, WL94);
sram_cell_6t_3 inst_cell_94_80 ( BL80, BLN80, WL94);
sram_cell_6t_3 inst_cell_94_79 ( BL79, BLN79, WL94);
sram_cell_6t_3 inst_cell_94_78 ( BL78, BLN78, WL94);
sram_cell_6t_3 inst_cell_94_77 ( BL77, BLN77, WL94);
sram_cell_6t_3 inst_cell_94_76 ( BL76, BLN76, WL94);
sram_cell_6t_3 inst_cell_94_75 ( BL75, BLN75, WL94);
sram_cell_6t_3 inst_cell_94_74 ( BL74, BLN74, WL94);
sram_cell_6t_3 inst_cell_94_73 ( BL73, BLN73, WL94);
sram_cell_6t_3 inst_cell_94_72 ( BL72, BLN72, WL94);
sram_cell_6t_3 inst_cell_94_71 ( BL71, BLN71, WL94);
sram_cell_6t_3 inst_cell_94_70 ( BL70, BLN70, WL94);
sram_cell_6t_3 inst_cell_94_69 ( BL69, BLN69, WL94);
sram_cell_6t_3 inst_cell_94_68 ( BL68, BLN68, WL94);
sram_cell_6t_3 inst_cell_94_67 ( BL67, BLN67, WL94);
sram_cell_6t_3 inst_cell_94_66 ( BL66, BLN66, WL94);
sram_cell_6t_3 inst_cell_94_65 ( BL65, BLN65, WL94);
sram_cell_6t_3 inst_cell_94_64 ( BL64, BLN64, WL94);
sram_cell_6t_3 inst_cell_94_63 ( BL63, BLN63, WL94);
sram_cell_6t_3 inst_cell_94_62 ( BL62, BLN62, WL94);
sram_cell_6t_3 inst_cell_94_61 ( BL61, BLN61, WL94);
sram_cell_6t_3 inst_cell_94_60 ( BL60, BLN60, WL94);
sram_cell_6t_3 inst_cell_94_59 ( BL59, BLN59, WL94);
sram_cell_6t_3 inst_cell_94_58 ( BL58, BLN58, WL94);
sram_cell_6t_3 inst_cell_94_57 ( BL57, BLN57, WL94);
sram_cell_6t_3 inst_cell_94_56 ( BL56, BLN56, WL94);
sram_cell_6t_3 inst_cell_94_55 ( BL55, BLN55, WL94);
sram_cell_6t_3 inst_cell_94_54 ( BL54, BLN54, WL94);
sram_cell_6t_3 inst_cell_94_53 ( BL53, BLN53, WL94);
sram_cell_6t_3 inst_cell_94_52 ( BL52, BLN52, WL94);
sram_cell_6t_3 inst_cell_94_51 ( BL51, BLN51, WL94);
sram_cell_6t_3 inst_cell_94_50 ( BL50, BLN50, WL94);
sram_cell_6t_3 inst_cell_94_49 ( BL49, BLN49, WL94);
sram_cell_6t_3 inst_cell_94_48 ( BL48, BLN48, WL94);
sram_cell_6t_3 inst_cell_94_47 ( BL47, BLN47, WL94);
sram_cell_6t_3 inst_cell_94_46 ( BL46, BLN46, WL94);
sram_cell_6t_3 inst_cell_94_45 ( BL45, BLN45, WL94);
sram_cell_6t_3 inst_cell_94_44 ( BL44, BLN44, WL94);
sram_cell_6t_3 inst_cell_94_43 ( BL43, BLN43, WL94);
sram_cell_6t_3 inst_cell_94_42 ( BL42, BLN42, WL94);
sram_cell_6t_3 inst_cell_94_41 ( BL41, BLN41, WL94);
sram_cell_6t_3 inst_cell_94_40 ( BL40, BLN40, WL94);
sram_cell_6t_3 inst_cell_94_39 ( BL39, BLN39, WL94);
sram_cell_6t_3 inst_cell_94_38 ( BL38, BLN38, WL94);
sram_cell_6t_3 inst_cell_94_37 ( BL37, BLN37, WL94);
sram_cell_6t_3 inst_cell_94_36 ( BL36, BLN36, WL94);
sram_cell_6t_3 inst_cell_94_35 ( BL35, BLN35, WL94);
sram_cell_6t_3 inst_cell_94_34 ( BL34, BLN34, WL94);
sram_cell_6t_3 inst_cell_94_33 ( BL33, BLN33, WL94);
sram_cell_6t_3 inst_cell_94_32 ( BL32, BLN32, WL94);
sram_cell_6t_3 inst_cell_94_31 ( BL31, BLN31, WL94);
sram_cell_6t_3 inst_cell_94_30 ( BL30, BLN30, WL94);
sram_cell_6t_3 inst_cell_94_29 ( BL29, BLN29, WL94);
sram_cell_6t_3 inst_cell_94_28 ( BL28, BLN28, WL94);
sram_cell_6t_3 inst_cell_94_27 ( BL27, BLN27, WL94);
sram_cell_6t_3 inst_cell_94_26 ( BL26, BLN26, WL94);
sram_cell_6t_3 inst_cell_94_25 ( BL25, BLN25, WL94);
sram_cell_6t_3 inst_cell_94_24 ( BL24, BLN24, WL94);
sram_cell_6t_3 inst_cell_94_23 ( BL23, BLN23, WL94);
sram_cell_6t_3 inst_cell_94_22 ( BL22, BLN22, WL94);
sram_cell_6t_3 inst_cell_94_21 ( BL21, BLN21, WL94);
sram_cell_6t_3 inst_cell_94_20 ( BL20, BLN20, WL94);
sram_cell_6t_3 inst_cell_94_19 ( BL19, BLN19, WL94);
sram_cell_6t_3 inst_cell_94_18 ( BL18, BLN18, WL94);
sram_cell_6t_3 inst_cell_94_17 ( BL17, BLN17, WL94);
sram_cell_6t_3 inst_cell_94_16 ( BL16, BLN16, WL94);
sram_cell_6t_3 inst_cell_94_15 ( BL15, BLN15, WL94);
sram_cell_6t_3 inst_cell_94_14 ( BL14, BLN14, WL94);
sram_cell_6t_3 inst_cell_94_13 ( BL13, BLN13, WL94);
sram_cell_6t_3 inst_cell_94_12 ( BL12, BLN12, WL94);
sram_cell_6t_3 inst_cell_94_11 ( BL11, BLN11, WL94);
sram_cell_6t_3 inst_cell_94_10 ( BL10, BLN10, WL94);
sram_cell_6t_3 inst_cell_94_9 ( BL9, BLN9, WL94);
sram_cell_6t_3 inst_cell_94_8 ( BL8, BLN8, WL94);
sram_cell_6t_3 inst_cell_94_7 ( BL7, BLN7, WL94);
sram_cell_6t_3 inst_cell_94_6 ( BL6, BLN6, WL94);
sram_cell_6t_3 inst_cell_94_5 ( BL5, BLN5, WL94);
sram_cell_6t_3 inst_cell_94_4 ( BL4, BLN4, WL94);
sram_cell_6t_3 inst_cell_94_3 ( BL3, BLN3, WL94);
sram_cell_6t_3 inst_cell_94_2 ( BL2, BLN2, WL94);
sram_cell_6t_3 inst_cell_94_1 ( BL1, BLN1, WL94);
sram_cell_6t_3 inst_cell_94_0 ( BL0, BLN0, WL94);
sram_cell_6t_3 inst_cell_93_127 ( BL127, BLN127, WL93);
sram_cell_6t_3 inst_cell_93_126 ( BL126, BLN126, WL93);
sram_cell_6t_3 inst_cell_93_125 ( BL125, BLN125, WL93);
sram_cell_6t_3 inst_cell_93_124 ( BL124, BLN124, WL93);
sram_cell_6t_3 inst_cell_93_123 ( BL123, BLN123, WL93);
sram_cell_6t_3 inst_cell_93_122 ( BL122, BLN122, WL93);
sram_cell_6t_3 inst_cell_93_121 ( BL121, BLN121, WL93);
sram_cell_6t_3 inst_cell_93_120 ( BL120, BLN120, WL93);
sram_cell_6t_3 inst_cell_93_119 ( BL119, BLN119, WL93);
sram_cell_6t_3 inst_cell_93_118 ( BL118, BLN118, WL93);
sram_cell_6t_3 inst_cell_93_117 ( BL117, BLN117, WL93);
sram_cell_6t_3 inst_cell_93_116 ( BL116, BLN116, WL93);
sram_cell_6t_3 inst_cell_93_115 ( BL115, BLN115, WL93);
sram_cell_6t_3 inst_cell_93_114 ( BL114, BLN114, WL93);
sram_cell_6t_3 inst_cell_93_113 ( BL113, BLN113, WL93);
sram_cell_6t_3 inst_cell_93_112 ( BL112, BLN112, WL93);
sram_cell_6t_3 inst_cell_93_111 ( BL111, BLN111, WL93);
sram_cell_6t_3 inst_cell_93_110 ( BL110, BLN110, WL93);
sram_cell_6t_3 inst_cell_93_109 ( BL109, BLN109, WL93);
sram_cell_6t_3 inst_cell_93_108 ( BL108, BLN108, WL93);
sram_cell_6t_3 inst_cell_93_107 ( BL107, BLN107, WL93);
sram_cell_6t_3 inst_cell_93_106 ( BL106, BLN106, WL93);
sram_cell_6t_3 inst_cell_93_105 ( BL105, BLN105, WL93);
sram_cell_6t_3 inst_cell_93_104 ( BL104, BLN104, WL93);
sram_cell_6t_3 inst_cell_93_103 ( BL103, BLN103, WL93);
sram_cell_6t_3 inst_cell_93_102 ( BL102, BLN102, WL93);
sram_cell_6t_3 inst_cell_93_101 ( BL101, BLN101, WL93);
sram_cell_6t_3 inst_cell_93_100 ( BL100, BLN100, WL93);
sram_cell_6t_3 inst_cell_93_99 ( BL99, BLN99, WL93);
sram_cell_6t_3 inst_cell_93_98 ( BL98, BLN98, WL93);
sram_cell_6t_3 inst_cell_93_97 ( BL97, BLN97, WL93);
sram_cell_6t_3 inst_cell_93_96 ( BL96, BLN96, WL93);
sram_cell_6t_3 inst_cell_93_95 ( BL95, BLN95, WL93);
sram_cell_6t_3 inst_cell_93_94 ( BL94, BLN94, WL93);
sram_cell_6t_3 inst_cell_93_93 ( BL93, BLN93, WL93);
sram_cell_6t_3 inst_cell_93_92 ( BL92, BLN92, WL93);
sram_cell_6t_3 inst_cell_93_91 ( BL91, BLN91, WL93);
sram_cell_6t_3 inst_cell_93_90 ( BL90, BLN90, WL93);
sram_cell_6t_3 inst_cell_93_89 ( BL89, BLN89, WL93);
sram_cell_6t_3 inst_cell_93_88 ( BL88, BLN88, WL93);
sram_cell_6t_3 inst_cell_93_87 ( BL87, BLN87, WL93);
sram_cell_6t_3 inst_cell_93_86 ( BL86, BLN86, WL93);
sram_cell_6t_3 inst_cell_93_85 ( BL85, BLN85, WL93);
sram_cell_6t_3 inst_cell_93_84 ( BL84, BLN84, WL93);
sram_cell_6t_3 inst_cell_93_83 ( BL83, BLN83, WL93);
sram_cell_6t_3 inst_cell_93_82 ( BL82, BLN82, WL93);
sram_cell_6t_3 inst_cell_93_81 ( BL81, BLN81, WL93);
sram_cell_6t_3 inst_cell_93_80 ( BL80, BLN80, WL93);
sram_cell_6t_3 inst_cell_93_79 ( BL79, BLN79, WL93);
sram_cell_6t_3 inst_cell_93_78 ( BL78, BLN78, WL93);
sram_cell_6t_3 inst_cell_93_77 ( BL77, BLN77, WL93);
sram_cell_6t_3 inst_cell_93_76 ( BL76, BLN76, WL93);
sram_cell_6t_3 inst_cell_93_75 ( BL75, BLN75, WL93);
sram_cell_6t_3 inst_cell_93_74 ( BL74, BLN74, WL93);
sram_cell_6t_3 inst_cell_93_73 ( BL73, BLN73, WL93);
sram_cell_6t_3 inst_cell_93_72 ( BL72, BLN72, WL93);
sram_cell_6t_3 inst_cell_93_71 ( BL71, BLN71, WL93);
sram_cell_6t_3 inst_cell_93_70 ( BL70, BLN70, WL93);
sram_cell_6t_3 inst_cell_93_69 ( BL69, BLN69, WL93);
sram_cell_6t_3 inst_cell_93_68 ( BL68, BLN68, WL93);
sram_cell_6t_3 inst_cell_93_67 ( BL67, BLN67, WL93);
sram_cell_6t_3 inst_cell_93_66 ( BL66, BLN66, WL93);
sram_cell_6t_3 inst_cell_93_65 ( BL65, BLN65, WL93);
sram_cell_6t_3 inst_cell_93_64 ( BL64, BLN64, WL93);
sram_cell_6t_3 inst_cell_93_63 ( BL63, BLN63, WL93);
sram_cell_6t_3 inst_cell_93_62 ( BL62, BLN62, WL93);
sram_cell_6t_3 inst_cell_93_61 ( BL61, BLN61, WL93);
sram_cell_6t_3 inst_cell_93_60 ( BL60, BLN60, WL93);
sram_cell_6t_3 inst_cell_93_59 ( BL59, BLN59, WL93);
sram_cell_6t_3 inst_cell_93_58 ( BL58, BLN58, WL93);
sram_cell_6t_3 inst_cell_93_57 ( BL57, BLN57, WL93);
sram_cell_6t_3 inst_cell_93_56 ( BL56, BLN56, WL93);
sram_cell_6t_3 inst_cell_93_55 ( BL55, BLN55, WL93);
sram_cell_6t_3 inst_cell_93_54 ( BL54, BLN54, WL93);
sram_cell_6t_3 inst_cell_93_53 ( BL53, BLN53, WL93);
sram_cell_6t_3 inst_cell_93_52 ( BL52, BLN52, WL93);
sram_cell_6t_3 inst_cell_93_51 ( BL51, BLN51, WL93);
sram_cell_6t_3 inst_cell_93_50 ( BL50, BLN50, WL93);
sram_cell_6t_3 inst_cell_93_49 ( BL49, BLN49, WL93);
sram_cell_6t_3 inst_cell_93_48 ( BL48, BLN48, WL93);
sram_cell_6t_3 inst_cell_93_47 ( BL47, BLN47, WL93);
sram_cell_6t_3 inst_cell_93_46 ( BL46, BLN46, WL93);
sram_cell_6t_3 inst_cell_93_45 ( BL45, BLN45, WL93);
sram_cell_6t_3 inst_cell_93_44 ( BL44, BLN44, WL93);
sram_cell_6t_3 inst_cell_93_43 ( BL43, BLN43, WL93);
sram_cell_6t_3 inst_cell_93_42 ( BL42, BLN42, WL93);
sram_cell_6t_3 inst_cell_93_41 ( BL41, BLN41, WL93);
sram_cell_6t_3 inst_cell_93_40 ( BL40, BLN40, WL93);
sram_cell_6t_3 inst_cell_93_39 ( BL39, BLN39, WL93);
sram_cell_6t_3 inst_cell_93_38 ( BL38, BLN38, WL93);
sram_cell_6t_3 inst_cell_93_37 ( BL37, BLN37, WL93);
sram_cell_6t_3 inst_cell_93_36 ( BL36, BLN36, WL93);
sram_cell_6t_3 inst_cell_93_35 ( BL35, BLN35, WL93);
sram_cell_6t_3 inst_cell_93_34 ( BL34, BLN34, WL93);
sram_cell_6t_3 inst_cell_93_33 ( BL33, BLN33, WL93);
sram_cell_6t_3 inst_cell_93_32 ( BL32, BLN32, WL93);
sram_cell_6t_3 inst_cell_93_31 ( BL31, BLN31, WL93);
sram_cell_6t_3 inst_cell_93_30 ( BL30, BLN30, WL93);
sram_cell_6t_3 inst_cell_93_29 ( BL29, BLN29, WL93);
sram_cell_6t_3 inst_cell_93_28 ( BL28, BLN28, WL93);
sram_cell_6t_3 inst_cell_93_27 ( BL27, BLN27, WL93);
sram_cell_6t_3 inst_cell_93_26 ( BL26, BLN26, WL93);
sram_cell_6t_3 inst_cell_93_25 ( BL25, BLN25, WL93);
sram_cell_6t_3 inst_cell_93_24 ( BL24, BLN24, WL93);
sram_cell_6t_3 inst_cell_93_23 ( BL23, BLN23, WL93);
sram_cell_6t_3 inst_cell_93_22 ( BL22, BLN22, WL93);
sram_cell_6t_3 inst_cell_93_21 ( BL21, BLN21, WL93);
sram_cell_6t_3 inst_cell_93_20 ( BL20, BLN20, WL93);
sram_cell_6t_3 inst_cell_93_19 ( BL19, BLN19, WL93);
sram_cell_6t_3 inst_cell_93_18 ( BL18, BLN18, WL93);
sram_cell_6t_3 inst_cell_93_17 ( BL17, BLN17, WL93);
sram_cell_6t_3 inst_cell_93_16 ( BL16, BLN16, WL93);
sram_cell_6t_3 inst_cell_93_15 ( BL15, BLN15, WL93);
sram_cell_6t_3 inst_cell_93_14 ( BL14, BLN14, WL93);
sram_cell_6t_3 inst_cell_93_13 ( BL13, BLN13, WL93);
sram_cell_6t_3 inst_cell_93_12 ( BL12, BLN12, WL93);
sram_cell_6t_3 inst_cell_93_11 ( BL11, BLN11, WL93);
sram_cell_6t_3 inst_cell_93_10 ( BL10, BLN10, WL93);
sram_cell_6t_3 inst_cell_93_9 ( BL9, BLN9, WL93);
sram_cell_6t_3 inst_cell_93_8 ( BL8, BLN8, WL93);
sram_cell_6t_3 inst_cell_93_7 ( BL7, BLN7, WL93);
sram_cell_6t_3 inst_cell_93_6 ( BL6, BLN6, WL93);
sram_cell_6t_3 inst_cell_93_5 ( BL5, BLN5, WL93);
sram_cell_6t_3 inst_cell_93_4 ( BL4, BLN4, WL93);
sram_cell_6t_3 inst_cell_93_3 ( BL3, BLN3, WL93);
sram_cell_6t_3 inst_cell_93_2 ( BL2, BLN2, WL93);
sram_cell_6t_3 inst_cell_93_1 ( BL1, BLN1, WL93);
sram_cell_6t_3 inst_cell_93_0 ( BL0, BLN0, WL93);
sram_cell_6t_3 inst_cell_92_127 ( BL127, BLN127, WL92);
sram_cell_6t_3 inst_cell_92_126 ( BL126, BLN126, WL92);
sram_cell_6t_3 inst_cell_92_125 ( BL125, BLN125, WL92);
sram_cell_6t_3 inst_cell_92_124 ( BL124, BLN124, WL92);
sram_cell_6t_3 inst_cell_92_123 ( BL123, BLN123, WL92);
sram_cell_6t_3 inst_cell_92_122 ( BL122, BLN122, WL92);
sram_cell_6t_3 inst_cell_92_121 ( BL121, BLN121, WL92);
sram_cell_6t_3 inst_cell_92_120 ( BL120, BLN120, WL92);
sram_cell_6t_3 inst_cell_92_119 ( BL119, BLN119, WL92);
sram_cell_6t_3 inst_cell_92_118 ( BL118, BLN118, WL92);
sram_cell_6t_3 inst_cell_92_117 ( BL117, BLN117, WL92);
sram_cell_6t_3 inst_cell_92_116 ( BL116, BLN116, WL92);
sram_cell_6t_3 inst_cell_92_115 ( BL115, BLN115, WL92);
sram_cell_6t_3 inst_cell_92_114 ( BL114, BLN114, WL92);
sram_cell_6t_3 inst_cell_92_113 ( BL113, BLN113, WL92);
sram_cell_6t_3 inst_cell_92_112 ( BL112, BLN112, WL92);
sram_cell_6t_3 inst_cell_92_111 ( BL111, BLN111, WL92);
sram_cell_6t_3 inst_cell_92_110 ( BL110, BLN110, WL92);
sram_cell_6t_3 inst_cell_92_109 ( BL109, BLN109, WL92);
sram_cell_6t_3 inst_cell_92_108 ( BL108, BLN108, WL92);
sram_cell_6t_3 inst_cell_92_107 ( BL107, BLN107, WL92);
sram_cell_6t_3 inst_cell_92_106 ( BL106, BLN106, WL92);
sram_cell_6t_3 inst_cell_92_105 ( BL105, BLN105, WL92);
sram_cell_6t_3 inst_cell_92_104 ( BL104, BLN104, WL92);
sram_cell_6t_3 inst_cell_92_103 ( BL103, BLN103, WL92);
sram_cell_6t_3 inst_cell_92_102 ( BL102, BLN102, WL92);
sram_cell_6t_3 inst_cell_92_101 ( BL101, BLN101, WL92);
sram_cell_6t_3 inst_cell_92_100 ( BL100, BLN100, WL92);
sram_cell_6t_3 inst_cell_92_99 ( BL99, BLN99, WL92);
sram_cell_6t_3 inst_cell_92_98 ( BL98, BLN98, WL92);
sram_cell_6t_3 inst_cell_92_97 ( BL97, BLN97, WL92);
sram_cell_6t_3 inst_cell_92_96 ( BL96, BLN96, WL92);
sram_cell_6t_3 inst_cell_92_95 ( BL95, BLN95, WL92);
sram_cell_6t_3 inst_cell_92_94 ( BL94, BLN94, WL92);
sram_cell_6t_3 inst_cell_92_93 ( BL93, BLN93, WL92);
sram_cell_6t_3 inst_cell_92_92 ( BL92, BLN92, WL92);
sram_cell_6t_3 inst_cell_92_91 ( BL91, BLN91, WL92);
sram_cell_6t_3 inst_cell_92_90 ( BL90, BLN90, WL92);
sram_cell_6t_3 inst_cell_92_89 ( BL89, BLN89, WL92);
sram_cell_6t_3 inst_cell_92_88 ( BL88, BLN88, WL92);
sram_cell_6t_3 inst_cell_92_87 ( BL87, BLN87, WL92);
sram_cell_6t_3 inst_cell_92_86 ( BL86, BLN86, WL92);
sram_cell_6t_3 inst_cell_92_85 ( BL85, BLN85, WL92);
sram_cell_6t_3 inst_cell_92_84 ( BL84, BLN84, WL92);
sram_cell_6t_3 inst_cell_92_83 ( BL83, BLN83, WL92);
sram_cell_6t_3 inst_cell_92_82 ( BL82, BLN82, WL92);
sram_cell_6t_3 inst_cell_92_81 ( BL81, BLN81, WL92);
sram_cell_6t_3 inst_cell_92_80 ( BL80, BLN80, WL92);
sram_cell_6t_3 inst_cell_92_79 ( BL79, BLN79, WL92);
sram_cell_6t_3 inst_cell_92_78 ( BL78, BLN78, WL92);
sram_cell_6t_3 inst_cell_92_77 ( BL77, BLN77, WL92);
sram_cell_6t_3 inst_cell_92_76 ( BL76, BLN76, WL92);
sram_cell_6t_3 inst_cell_92_75 ( BL75, BLN75, WL92);
sram_cell_6t_3 inst_cell_92_74 ( BL74, BLN74, WL92);
sram_cell_6t_3 inst_cell_92_73 ( BL73, BLN73, WL92);
sram_cell_6t_3 inst_cell_92_72 ( BL72, BLN72, WL92);
sram_cell_6t_3 inst_cell_92_71 ( BL71, BLN71, WL92);
sram_cell_6t_3 inst_cell_92_70 ( BL70, BLN70, WL92);
sram_cell_6t_3 inst_cell_92_69 ( BL69, BLN69, WL92);
sram_cell_6t_3 inst_cell_92_68 ( BL68, BLN68, WL92);
sram_cell_6t_3 inst_cell_92_67 ( BL67, BLN67, WL92);
sram_cell_6t_3 inst_cell_92_66 ( BL66, BLN66, WL92);
sram_cell_6t_3 inst_cell_92_65 ( BL65, BLN65, WL92);
sram_cell_6t_3 inst_cell_92_64 ( BL64, BLN64, WL92);
sram_cell_6t_3 inst_cell_92_63 ( BL63, BLN63, WL92);
sram_cell_6t_3 inst_cell_92_62 ( BL62, BLN62, WL92);
sram_cell_6t_3 inst_cell_92_61 ( BL61, BLN61, WL92);
sram_cell_6t_3 inst_cell_92_60 ( BL60, BLN60, WL92);
sram_cell_6t_3 inst_cell_92_59 ( BL59, BLN59, WL92);
sram_cell_6t_3 inst_cell_92_58 ( BL58, BLN58, WL92);
sram_cell_6t_3 inst_cell_92_57 ( BL57, BLN57, WL92);
sram_cell_6t_3 inst_cell_92_56 ( BL56, BLN56, WL92);
sram_cell_6t_3 inst_cell_92_55 ( BL55, BLN55, WL92);
sram_cell_6t_3 inst_cell_92_54 ( BL54, BLN54, WL92);
sram_cell_6t_3 inst_cell_92_53 ( BL53, BLN53, WL92);
sram_cell_6t_3 inst_cell_92_52 ( BL52, BLN52, WL92);
sram_cell_6t_3 inst_cell_92_51 ( BL51, BLN51, WL92);
sram_cell_6t_3 inst_cell_92_50 ( BL50, BLN50, WL92);
sram_cell_6t_3 inst_cell_92_49 ( BL49, BLN49, WL92);
sram_cell_6t_3 inst_cell_92_48 ( BL48, BLN48, WL92);
sram_cell_6t_3 inst_cell_92_47 ( BL47, BLN47, WL92);
sram_cell_6t_3 inst_cell_92_46 ( BL46, BLN46, WL92);
sram_cell_6t_3 inst_cell_92_45 ( BL45, BLN45, WL92);
sram_cell_6t_3 inst_cell_92_44 ( BL44, BLN44, WL92);
sram_cell_6t_3 inst_cell_92_43 ( BL43, BLN43, WL92);
sram_cell_6t_3 inst_cell_92_42 ( BL42, BLN42, WL92);
sram_cell_6t_3 inst_cell_92_41 ( BL41, BLN41, WL92);
sram_cell_6t_3 inst_cell_92_40 ( BL40, BLN40, WL92);
sram_cell_6t_3 inst_cell_92_39 ( BL39, BLN39, WL92);
sram_cell_6t_3 inst_cell_92_38 ( BL38, BLN38, WL92);
sram_cell_6t_3 inst_cell_92_37 ( BL37, BLN37, WL92);
sram_cell_6t_3 inst_cell_92_36 ( BL36, BLN36, WL92);
sram_cell_6t_3 inst_cell_92_35 ( BL35, BLN35, WL92);
sram_cell_6t_3 inst_cell_92_34 ( BL34, BLN34, WL92);
sram_cell_6t_3 inst_cell_92_33 ( BL33, BLN33, WL92);
sram_cell_6t_3 inst_cell_92_32 ( BL32, BLN32, WL92);
sram_cell_6t_3 inst_cell_92_31 ( BL31, BLN31, WL92);
sram_cell_6t_3 inst_cell_92_30 ( BL30, BLN30, WL92);
sram_cell_6t_3 inst_cell_92_29 ( BL29, BLN29, WL92);
sram_cell_6t_3 inst_cell_92_28 ( BL28, BLN28, WL92);
sram_cell_6t_3 inst_cell_92_27 ( BL27, BLN27, WL92);
sram_cell_6t_3 inst_cell_92_26 ( BL26, BLN26, WL92);
sram_cell_6t_3 inst_cell_92_25 ( BL25, BLN25, WL92);
sram_cell_6t_3 inst_cell_92_24 ( BL24, BLN24, WL92);
sram_cell_6t_3 inst_cell_92_23 ( BL23, BLN23, WL92);
sram_cell_6t_3 inst_cell_92_22 ( BL22, BLN22, WL92);
sram_cell_6t_3 inst_cell_92_21 ( BL21, BLN21, WL92);
sram_cell_6t_3 inst_cell_92_20 ( BL20, BLN20, WL92);
sram_cell_6t_3 inst_cell_92_19 ( BL19, BLN19, WL92);
sram_cell_6t_3 inst_cell_92_18 ( BL18, BLN18, WL92);
sram_cell_6t_3 inst_cell_92_17 ( BL17, BLN17, WL92);
sram_cell_6t_3 inst_cell_92_16 ( BL16, BLN16, WL92);
sram_cell_6t_3 inst_cell_92_15 ( BL15, BLN15, WL92);
sram_cell_6t_3 inst_cell_92_14 ( BL14, BLN14, WL92);
sram_cell_6t_3 inst_cell_92_13 ( BL13, BLN13, WL92);
sram_cell_6t_3 inst_cell_92_12 ( BL12, BLN12, WL92);
sram_cell_6t_3 inst_cell_92_11 ( BL11, BLN11, WL92);
sram_cell_6t_3 inst_cell_92_10 ( BL10, BLN10, WL92);
sram_cell_6t_3 inst_cell_92_9 ( BL9, BLN9, WL92);
sram_cell_6t_3 inst_cell_92_8 ( BL8, BLN8, WL92);
sram_cell_6t_3 inst_cell_92_7 ( BL7, BLN7, WL92);
sram_cell_6t_3 inst_cell_92_6 ( BL6, BLN6, WL92);
sram_cell_6t_3 inst_cell_92_5 ( BL5, BLN5, WL92);
sram_cell_6t_3 inst_cell_92_4 ( BL4, BLN4, WL92);
sram_cell_6t_3 inst_cell_92_3 ( BL3, BLN3, WL92);
sram_cell_6t_3 inst_cell_92_2 ( BL2, BLN2, WL92);
sram_cell_6t_3 inst_cell_92_1 ( BL1, BLN1, WL92);
sram_cell_6t_3 inst_cell_92_0 ( BL0, BLN0, WL92);
sram_cell_6t_3 inst_cell_91_127 ( BL127, BLN127, WL91);
sram_cell_6t_3 inst_cell_91_126 ( BL126, BLN126, WL91);
sram_cell_6t_3 inst_cell_91_125 ( BL125, BLN125, WL91);
sram_cell_6t_3 inst_cell_91_124 ( BL124, BLN124, WL91);
sram_cell_6t_3 inst_cell_91_123 ( BL123, BLN123, WL91);
sram_cell_6t_3 inst_cell_91_122 ( BL122, BLN122, WL91);
sram_cell_6t_3 inst_cell_91_121 ( BL121, BLN121, WL91);
sram_cell_6t_3 inst_cell_91_120 ( BL120, BLN120, WL91);
sram_cell_6t_3 inst_cell_91_119 ( BL119, BLN119, WL91);
sram_cell_6t_3 inst_cell_91_118 ( BL118, BLN118, WL91);
sram_cell_6t_3 inst_cell_91_117 ( BL117, BLN117, WL91);
sram_cell_6t_3 inst_cell_91_116 ( BL116, BLN116, WL91);
sram_cell_6t_3 inst_cell_91_115 ( BL115, BLN115, WL91);
sram_cell_6t_3 inst_cell_91_114 ( BL114, BLN114, WL91);
sram_cell_6t_3 inst_cell_91_113 ( BL113, BLN113, WL91);
sram_cell_6t_3 inst_cell_91_112 ( BL112, BLN112, WL91);
sram_cell_6t_3 inst_cell_91_111 ( BL111, BLN111, WL91);
sram_cell_6t_3 inst_cell_91_110 ( BL110, BLN110, WL91);
sram_cell_6t_3 inst_cell_91_109 ( BL109, BLN109, WL91);
sram_cell_6t_3 inst_cell_91_108 ( BL108, BLN108, WL91);
sram_cell_6t_3 inst_cell_91_107 ( BL107, BLN107, WL91);
sram_cell_6t_3 inst_cell_91_106 ( BL106, BLN106, WL91);
sram_cell_6t_3 inst_cell_91_105 ( BL105, BLN105, WL91);
sram_cell_6t_3 inst_cell_91_104 ( BL104, BLN104, WL91);
sram_cell_6t_3 inst_cell_91_103 ( BL103, BLN103, WL91);
sram_cell_6t_3 inst_cell_91_102 ( BL102, BLN102, WL91);
sram_cell_6t_3 inst_cell_91_101 ( BL101, BLN101, WL91);
sram_cell_6t_3 inst_cell_91_100 ( BL100, BLN100, WL91);
sram_cell_6t_3 inst_cell_91_99 ( BL99, BLN99, WL91);
sram_cell_6t_3 inst_cell_91_98 ( BL98, BLN98, WL91);
sram_cell_6t_3 inst_cell_91_97 ( BL97, BLN97, WL91);
sram_cell_6t_3 inst_cell_91_96 ( BL96, BLN96, WL91);
sram_cell_6t_3 inst_cell_91_95 ( BL95, BLN95, WL91);
sram_cell_6t_3 inst_cell_91_94 ( BL94, BLN94, WL91);
sram_cell_6t_3 inst_cell_91_93 ( BL93, BLN93, WL91);
sram_cell_6t_3 inst_cell_91_92 ( BL92, BLN92, WL91);
sram_cell_6t_3 inst_cell_91_91 ( BL91, BLN91, WL91);
sram_cell_6t_3 inst_cell_91_90 ( BL90, BLN90, WL91);
sram_cell_6t_3 inst_cell_91_89 ( BL89, BLN89, WL91);
sram_cell_6t_3 inst_cell_91_88 ( BL88, BLN88, WL91);
sram_cell_6t_3 inst_cell_91_87 ( BL87, BLN87, WL91);
sram_cell_6t_3 inst_cell_91_86 ( BL86, BLN86, WL91);
sram_cell_6t_3 inst_cell_91_85 ( BL85, BLN85, WL91);
sram_cell_6t_3 inst_cell_91_84 ( BL84, BLN84, WL91);
sram_cell_6t_3 inst_cell_91_83 ( BL83, BLN83, WL91);
sram_cell_6t_3 inst_cell_91_82 ( BL82, BLN82, WL91);
sram_cell_6t_3 inst_cell_91_81 ( BL81, BLN81, WL91);
sram_cell_6t_3 inst_cell_91_80 ( BL80, BLN80, WL91);
sram_cell_6t_3 inst_cell_91_79 ( BL79, BLN79, WL91);
sram_cell_6t_3 inst_cell_91_78 ( BL78, BLN78, WL91);
sram_cell_6t_3 inst_cell_91_77 ( BL77, BLN77, WL91);
sram_cell_6t_3 inst_cell_91_76 ( BL76, BLN76, WL91);
sram_cell_6t_3 inst_cell_91_75 ( BL75, BLN75, WL91);
sram_cell_6t_3 inst_cell_91_74 ( BL74, BLN74, WL91);
sram_cell_6t_3 inst_cell_91_73 ( BL73, BLN73, WL91);
sram_cell_6t_3 inst_cell_91_72 ( BL72, BLN72, WL91);
sram_cell_6t_3 inst_cell_91_71 ( BL71, BLN71, WL91);
sram_cell_6t_3 inst_cell_91_70 ( BL70, BLN70, WL91);
sram_cell_6t_3 inst_cell_91_69 ( BL69, BLN69, WL91);
sram_cell_6t_3 inst_cell_91_68 ( BL68, BLN68, WL91);
sram_cell_6t_3 inst_cell_91_67 ( BL67, BLN67, WL91);
sram_cell_6t_3 inst_cell_91_66 ( BL66, BLN66, WL91);
sram_cell_6t_3 inst_cell_91_65 ( BL65, BLN65, WL91);
sram_cell_6t_3 inst_cell_91_64 ( BL64, BLN64, WL91);
sram_cell_6t_3 inst_cell_91_63 ( BL63, BLN63, WL91);
sram_cell_6t_3 inst_cell_91_62 ( BL62, BLN62, WL91);
sram_cell_6t_3 inst_cell_91_61 ( BL61, BLN61, WL91);
sram_cell_6t_3 inst_cell_91_60 ( BL60, BLN60, WL91);
sram_cell_6t_3 inst_cell_91_59 ( BL59, BLN59, WL91);
sram_cell_6t_3 inst_cell_91_58 ( BL58, BLN58, WL91);
sram_cell_6t_3 inst_cell_91_57 ( BL57, BLN57, WL91);
sram_cell_6t_3 inst_cell_91_56 ( BL56, BLN56, WL91);
sram_cell_6t_3 inst_cell_91_55 ( BL55, BLN55, WL91);
sram_cell_6t_3 inst_cell_91_54 ( BL54, BLN54, WL91);
sram_cell_6t_3 inst_cell_91_53 ( BL53, BLN53, WL91);
sram_cell_6t_3 inst_cell_91_52 ( BL52, BLN52, WL91);
sram_cell_6t_3 inst_cell_91_51 ( BL51, BLN51, WL91);
sram_cell_6t_3 inst_cell_91_50 ( BL50, BLN50, WL91);
sram_cell_6t_3 inst_cell_91_49 ( BL49, BLN49, WL91);
sram_cell_6t_3 inst_cell_91_48 ( BL48, BLN48, WL91);
sram_cell_6t_3 inst_cell_91_47 ( BL47, BLN47, WL91);
sram_cell_6t_3 inst_cell_91_46 ( BL46, BLN46, WL91);
sram_cell_6t_3 inst_cell_91_45 ( BL45, BLN45, WL91);
sram_cell_6t_3 inst_cell_91_44 ( BL44, BLN44, WL91);
sram_cell_6t_3 inst_cell_91_43 ( BL43, BLN43, WL91);
sram_cell_6t_3 inst_cell_91_42 ( BL42, BLN42, WL91);
sram_cell_6t_3 inst_cell_91_41 ( BL41, BLN41, WL91);
sram_cell_6t_3 inst_cell_91_40 ( BL40, BLN40, WL91);
sram_cell_6t_3 inst_cell_91_39 ( BL39, BLN39, WL91);
sram_cell_6t_3 inst_cell_91_38 ( BL38, BLN38, WL91);
sram_cell_6t_3 inst_cell_91_37 ( BL37, BLN37, WL91);
sram_cell_6t_3 inst_cell_91_36 ( BL36, BLN36, WL91);
sram_cell_6t_3 inst_cell_91_35 ( BL35, BLN35, WL91);
sram_cell_6t_3 inst_cell_91_34 ( BL34, BLN34, WL91);
sram_cell_6t_3 inst_cell_91_33 ( BL33, BLN33, WL91);
sram_cell_6t_3 inst_cell_91_32 ( BL32, BLN32, WL91);
sram_cell_6t_3 inst_cell_91_31 ( BL31, BLN31, WL91);
sram_cell_6t_3 inst_cell_91_30 ( BL30, BLN30, WL91);
sram_cell_6t_3 inst_cell_91_29 ( BL29, BLN29, WL91);
sram_cell_6t_3 inst_cell_91_28 ( BL28, BLN28, WL91);
sram_cell_6t_3 inst_cell_91_27 ( BL27, BLN27, WL91);
sram_cell_6t_3 inst_cell_91_26 ( BL26, BLN26, WL91);
sram_cell_6t_3 inst_cell_91_25 ( BL25, BLN25, WL91);
sram_cell_6t_3 inst_cell_91_24 ( BL24, BLN24, WL91);
sram_cell_6t_3 inst_cell_91_23 ( BL23, BLN23, WL91);
sram_cell_6t_3 inst_cell_91_22 ( BL22, BLN22, WL91);
sram_cell_6t_3 inst_cell_91_21 ( BL21, BLN21, WL91);
sram_cell_6t_3 inst_cell_91_20 ( BL20, BLN20, WL91);
sram_cell_6t_3 inst_cell_91_19 ( BL19, BLN19, WL91);
sram_cell_6t_3 inst_cell_91_18 ( BL18, BLN18, WL91);
sram_cell_6t_3 inst_cell_91_17 ( BL17, BLN17, WL91);
sram_cell_6t_3 inst_cell_91_16 ( BL16, BLN16, WL91);
sram_cell_6t_3 inst_cell_91_15 ( BL15, BLN15, WL91);
sram_cell_6t_3 inst_cell_91_14 ( BL14, BLN14, WL91);
sram_cell_6t_3 inst_cell_91_13 ( BL13, BLN13, WL91);
sram_cell_6t_3 inst_cell_91_12 ( BL12, BLN12, WL91);
sram_cell_6t_3 inst_cell_91_11 ( BL11, BLN11, WL91);
sram_cell_6t_3 inst_cell_91_10 ( BL10, BLN10, WL91);
sram_cell_6t_3 inst_cell_91_9 ( BL9, BLN9, WL91);
sram_cell_6t_3 inst_cell_91_8 ( BL8, BLN8, WL91);
sram_cell_6t_3 inst_cell_91_7 ( BL7, BLN7, WL91);
sram_cell_6t_3 inst_cell_91_6 ( BL6, BLN6, WL91);
sram_cell_6t_3 inst_cell_91_5 ( BL5, BLN5, WL91);
sram_cell_6t_3 inst_cell_91_4 ( BL4, BLN4, WL91);
sram_cell_6t_3 inst_cell_91_3 ( BL3, BLN3, WL91);
sram_cell_6t_3 inst_cell_91_2 ( BL2, BLN2, WL91);
sram_cell_6t_3 inst_cell_91_1 ( BL1, BLN1, WL91);
sram_cell_6t_3 inst_cell_91_0 ( BL0, BLN0, WL91);
sram_cell_6t_3 inst_cell_90_127 ( BL127, BLN127, WL90);
sram_cell_6t_3 inst_cell_90_126 ( BL126, BLN126, WL90);
sram_cell_6t_3 inst_cell_90_125 ( BL125, BLN125, WL90);
sram_cell_6t_3 inst_cell_90_124 ( BL124, BLN124, WL90);
sram_cell_6t_3 inst_cell_90_123 ( BL123, BLN123, WL90);
sram_cell_6t_3 inst_cell_90_122 ( BL122, BLN122, WL90);
sram_cell_6t_3 inst_cell_90_121 ( BL121, BLN121, WL90);
sram_cell_6t_3 inst_cell_90_120 ( BL120, BLN120, WL90);
sram_cell_6t_3 inst_cell_90_119 ( BL119, BLN119, WL90);
sram_cell_6t_3 inst_cell_90_118 ( BL118, BLN118, WL90);
sram_cell_6t_3 inst_cell_90_117 ( BL117, BLN117, WL90);
sram_cell_6t_3 inst_cell_90_116 ( BL116, BLN116, WL90);
sram_cell_6t_3 inst_cell_90_115 ( BL115, BLN115, WL90);
sram_cell_6t_3 inst_cell_90_114 ( BL114, BLN114, WL90);
sram_cell_6t_3 inst_cell_90_113 ( BL113, BLN113, WL90);
sram_cell_6t_3 inst_cell_90_112 ( BL112, BLN112, WL90);
sram_cell_6t_3 inst_cell_90_111 ( BL111, BLN111, WL90);
sram_cell_6t_3 inst_cell_90_110 ( BL110, BLN110, WL90);
sram_cell_6t_3 inst_cell_90_109 ( BL109, BLN109, WL90);
sram_cell_6t_3 inst_cell_90_108 ( BL108, BLN108, WL90);
sram_cell_6t_3 inst_cell_90_107 ( BL107, BLN107, WL90);
sram_cell_6t_3 inst_cell_90_106 ( BL106, BLN106, WL90);
sram_cell_6t_3 inst_cell_90_105 ( BL105, BLN105, WL90);
sram_cell_6t_3 inst_cell_90_104 ( BL104, BLN104, WL90);
sram_cell_6t_3 inst_cell_90_103 ( BL103, BLN103, WL90);
sram_cell_6t_3 inst_cell_90_102 ( BL102, BLN102, WL90);
sram_cell_6t_3 inst_cell_90_101 ( BL101, BLN101, WL90);
sram_cell_6t_3 inst_cell_90_100 ( BL100, BLN100, WL90);
sram_cell_6t_3 inst_cell_90_99 ( BL99, BLN99, WL90);
sram_cell_6t_3 inst_cell_90_98 ( BL98, BLN98, WL90);
sram_cell_6t_3 inst_cell_90_97 ( BL97, BLN97, WL90);
sram_cell_6t_3 inst_cell_90_96 ( BL96, BLN96, WL90);
sram_cell_6t_3 inst_cell_90_95 ( BL95, BLN95, WL90);
sram_cell_6t_3 inst_cell_90_94 ( BL94, BLN94, WL90);
sram_cell_6t_3 inst_cell_90_93 ( BL93, BLN93, WL90);
sram_cell_6t_3 inst_cell_90_92 ( BL92, BLN92, WL90);
sram_cell_6t_3 inst_cell_90_91 ( BL91, BLN91, WL90);
sram_cell_6t_3 inst_cell_90_90 ( BL90, BLN90, WL90);
sram_cell_6t_3 inst_cell_90_89 ( BL89, BLN89, WL90);
sram_cell_6t_3 inst_cell_90_88 ( BL88, BLN88, WL90);
sram_cell_6t_3 inst_cell_90_87 ( BL87, BLN87, WL90);
sram_cell_6t_3 inst_cell_90_86 ( BL86, BLN86, WL90);
sram_cell_6t_3 inst_cell_90_85 ( BL85, BLN85, WL90);
sram_cell_6t_3 inst_cell_90_84 ( BL84, BLN84, WL90);
sram_cell_6t_3 inst_cell_90_83 ( BL83, BLN83, WL90);
sram_cell_6t_3 inst_cell_90_82 ( BL82, BLN82, WL90);
sram_cell_6t_3 inst_cell_90_81 ( BL81, BLN81, WL90);
sram_cell_6t_3 inst_cell_90_80 ( BL80, BLN80, WL90);
sram_cell_6t_3 inst_cell_90_79 ( BL79, BLN79, WL90);
sram_cell_6t_3 inst_cell_90_78 ( BL78, BLN78, WL90);
sram_cell_6t_3 inst_cell_90_77 ( BL77, BLN77, WL90);
sram_cell_6t_3 inst_cell_90_76 ( BL76, BLN76, WL90);
sram_cell_6t_3 inst_cell_90_75 ( BL75, BLN75, WL90);
sram_cell_6t_3 inst_cell_90_74 ( BL74, BLN74, WL90);
sram_cell_6t_3 inst_cell_90_73 ( BL73, BLN73, WL90);
sram_cell_6t_3 inst_cell_90_72 ( BL72, BLN72, WL90);
sram_cell_6t_3 inst_cell_90_71 ( BL71, BLN71, WL90);
sram_cell_6t_3 inst_cell_90_70 ( BL70, BLN70, WL90);
sram_cell_6t_3 inst_cell_90_69 ( BL69, BLN69, WL90);
sram_cell_6t_3 inst_cell_90_68 ( BL68, BLN68, WL90);
sram_cell_6t_3 inst_cell_90_67 ( BL67, BLN67, WL90);
sram_cell_6t_3 inst_cell_90_66 ( BL66, BLN66, WL90);
sram_cell_6t_3 inst_cell_90_65 ( BL65, BLN65, WL90);
sram_cell_6t_3 inst_cell_90_64 ( BL64, BLN64, WL90);
sram_cell_6t_3 inst_cell_90_63 ( BL63, BLN63, WL90);
sram_cell_6t_3 inst_cell_90_62 ( BL62, BLN62, WL90);
sram_cell_6t_3 inst_cell_90_61 ( BL61, BLN61, WL90);
sram_cell_6t_3 inst_cell_90_60 ( BL60, BLN60, WL90);
sram_cell_6t_3 inst_cell_90_59 ( BL59, BLN59, WL90);
sram_cell_6t_3 inst_cell_90_58 ( BL58, BLN58, WL90);
sram_cell_6t_3 inst_cell_90_57 ( BL57, BLN57, WL90);
sram_cell_6t_3 inst_cell_90_56 ( BL56, BLN56, WL90);
sram_cell_6t_3 inst_cell_90_55 ( BL55, BLN55, WL90);
sram_cell_6t_3 inst_cell_90_54 ( BL54, BLN54, WL90);
sram_cell_6t_3 inst_cell_90_53 ( BL53, BLN53, WL90);
sram_cell_6t_3 inst_cell_90_52 ( BL52, BLN52, WL90);
sram_cell_6t_3 inst_cell_90_51 ( BL51, BLN51, WL90);
sram_cell_6t_3 inst_cell_90_50 ( BL50, BLN50, WL90);
sram_cell_6t_3 inst_cell_90_49 ( BL49, BLN49, WL90);
sram_cell_6t_3 inst_cell_90_48 ( BL48, BLN48, WL90);
sram_cell_6t_3 inst_cell_90_47 ( BL47, BLN47, WL90);
sram_cell_6t_3 inst_cell_90_46 ( BL46, BLN46, WL90);
sram_cell_6t_3 inst_cell_90_45 ( BL45, BLN45, WL90);
sram_cell_6t_3 inst_cell_90_44 ( BL44, BLN44, WL90);
sram_cell_6t_3 inst_cell_90_43 ( BL43, BLN43, WL90);
sram_cell_6t_3 inst_cell_90_42 ( BL42, BLN42, WL90);
sram_cell_6t_3 inst_cell_90_41 ( BL41, BLN41, WL90);
sram_cell_6t_3 inst_cell_90_40 ( BL40, BLN40, WL90);
sram_cell_6t_3 inst_cell_90_39 ( BL39, BLN39, WL90);
sram_cell_6t_3 inst_cell_90_38 ( BL38, BLN38, WL90);
sram_cell_6t_3 inst_cell_90_37 ( BL37, BLN37, WL90);
sram_cell_6t_3 inst_cell_90_36 ( BL36, BLN36, WL90);
sram_cell_6t_3 inst_cell_90_35 ( BL35, BLN35, WL90);
sram_cell_6t_3 inst_cell_90_34 ( BL34, BLN34, WL90);
sram_cell_6t_3 inst_cell_90_33 ( BL33, BLN33, WL90);
sram_cell_6t_3 inst_cell_90_32 ( BL32, BLN32, WL90);
sram_cell_6t_3 inst_cell_90_31 ( BL31, BLN31, WL90);
sram_cell_6t_3 inst_cell_90_30 ( BL30, BLN30, WL90);
sram_cell_6t_3 inst_cell_90_29 ( BL29, BLN29, WL90);
sram_cell_6t_3 inst_cell_90_28 ( BL28, BLN28, WL90);
sram_cell_6t_3 inst_cell_90_27 ( BL27, BLN27, WL90);
sram_cell_6t_3 inst_cell_90_26 ( BL26, BLN26, WL90);
sram_cell_6t_3 inst_cell_90_25 ( BL25, BLN25, WL90);
sram_cell_6t_3 inst_cell_90_24 ( BL24, BLN24, WL90);
sram_cell_6t_3 inst_cell_90_23 ( BL23, BLN23, WL90);
sram_cell_6t_3 inst_cell_90_22 ( BL22, BLN22, WL90);
sram_cell_6t_3 inst_cell_90_21 ( BL21, BLN21, WL90);
sram_cell_6t_3 inst_cell_90_20 ( BL20, BLN20, WL90);
sram_cell_6t_3 inst_cell_90_19 ( BL19, BLN19, WL90);
sram_cell_6t_3 inst_cell_90_18 ( BL18, BLN18, WL90);
sram_cell_6t_3 inst_cell_90_17 ( BL17, BLN17, WL90);
sram_cell_6t_3 inst_cell_90_16 ( BL16, BLN16, WL90);
sram_cell_6t_3 inst_cell_90_15 ( BL15, BLN15, WL90);
sram_cell_6t_3 inst_cell_90_14 ( BL14, BLN14, WL90);
sram_cell_6t_3 inst_cell_90_13 ( BL13, BLN13, WL90);
sram_cell_6t_3 inst_cell_90_12 ( BL12, BLN12, WL90);
sram_cell_6t_3 inst_cell_90_11 ( BL11, BLN11, WL90);
sram_cell_6t_3 inst_cell_90_10 ( BL10, BLN10, WL90);
sram_cell_6t_3 inst_cell_90_9 ( BL9, BLN9, WL90);
sram_cell_6t_3 inst_cell_90_8 ( BL8, BLN8, WL90);
sram_cell_6t_3 inst_cell_90_7 ( BL7, BLN7, WL90);
sram_cell_6t_3 inst_cell_90_6 ( BL6, BLN6, WL90);
sram_cell_6t_3 inst_cell_90_5 ( BL5, BLN5, WL90);
sram_cell_6t_3 inst_cell_90_4 ( BL4, BLN4, WL90);
sram_cell_6t_3 inst_cell_90_3 ( BL3, BLN3, WL90);
sram_cell_6t_3 inst_cell_90_2 ( BL2, BLN2, WL90);
sram_cell_6t_3 inst_cell_90_1 ( BL1, BLN1, WL90);
sram_cell_6t_3 inst_cell_90_0 ( BL0, BLN0, WL90);
sram_cell_6t_3 inst_cell_89_127 ( BL127, BLN127, WL89);
sram_cell_6t_3 inst_cell_89_126 ( BL126, BLN126, WL89);
sram_cell_6t_3 inst_cell_89_125 ( BL125, BLN125, WL89);
sram_cell_6t_3 inst_cell_89_124 ( BL124, BLN124, WL89);
sram_cell_6t_3 inst_cell_89_123 ( BL123, BLN123, WL89);
sram_cell_6t_3 inst_cell_89_122 ( BL122, BLN122, WL89);
sram_cell_6t_3 inst_cell_89_121 ( BL121, BLN121, WL89);
sram_cell_6t_3 inst_cell_89_120 ( BL120, BLN120, WL89);
sram_cell_6t_3 inst_cell_89_119 ( BL119, BLN119, WL89);
sram_cell_6t_3 inst_cell_89_118 ( BL118, BLN118, WL89);
sram_cell_6t_3 inst_cell_89_117 ( BL117, BLN117, WL89);
sram_cell_6t_3 inst_cell_89_116 ( BL116, BLN116, WL89);
sram_cell_6t_3 inst_cell_89_115 ( BL115, BLN115, WL89);
sram_cell_6t_3 inst_cell_89_114 ( BL114, BLN114, WL89);
sram_cell_6t_3 inst_cell_89_113 ( BL113, BLN113, WL89);
sram_cell_6t_3 inst_cell_89_112 ( BL112, BLN112, WL89);
sram_cell_6t_3 inst_cell_89_111 ( BL111, BLN111, WL89);
sram_cell_6t_3 inst_cell_89_110 ( BL110, BLN110, WL89);
sram_cell_6t_3 inst_cell_89_109 ( BL109, BLN109, WL89);
sram_cell_6t_3 inst_cell_89_108 ( BL108, BLN108, WL89);
sram_cell_6t_3 inst_cell_89_107 ( BL107, BLN107, WL89);
sram_cell_6t_3 inst_cell_89_106 ( BL106, BLN106, WL89);
sram_cell_6t_3 inst_cell_89_105 ( BL105, BLN105, WL89);
sram_cell_6t_3 inst_cell_89_104 ( BL104, BLN104, WL89);
sram_cell_6t_3 inst_cell_89_103 ( BL103, BLN103, WL89);
sram_cell_6t_3 inst_cell_89_102 ( BL102, BLN102, WL89);
sram_cell_6t_3 inst_cell_89_101 ( BL101, BLN101, WL89);
sram_cell_6t_3 inst_cell_89_100 ( BL100, BLN100, WL89);
sram_cell_6t_3 inst_cell_89_99 ( BL99, BLN99, WL89);
sram_cell_6t_3 inst_cell_89_98 ( BL98, BLN98, WL89);
sram_cell_6t_3 inst_cell_89_97 ( BL97, BLN97, WL89);
sram_cell_6t_3 inst_cell_89_96 ( BL96, BLN96, WL89);
sram_cell_6t_3 inst_cell_89_95 ( BL95, BLN95, WL89);
sram_cell_6t_3 inst_cell_89_94 ( BL94, BLN94, WL89);
sram_cell_6t_3 inst_cell_89_93 ( BL93, BLN93, WL89);
sram_cell_6t_3 inst_cell_89_92 ( BL92, BLN92, WL89);
sram_cell_6t_3 inst_cell_89_91 ( BL91, BLN91, WL89);
sram_cell_6t_3 inst_cell_89_90 ( BL90, BLN90, WL89);
sram_cell_6t_3 inst_cell_89_89 ( BL89, BLN89, WL89);
sram_cell_6t_3 inst_cell_89_88 ( BL88, BLN88, WL89);
sram_cell_6t_3 inst_cell_89_87 ( BL87, BLN87, WL89);
sram_cell_6t_3 inst_cell_89_86 ( BL86, BLN86, WL89);
sram_cell_6t_3 inst_cell_89_85 ( BL85, BLN85, WL89);
sram_cell_6t_3 inst_cell_89_84 ( BL84, BLN84, WL89);
sram_cell_6t_3 inst_cell_89_83 ( BL83, BLN83, WL89);
sram_cell_6t_3 inst_cell_89_82 ( BL82, BLN82, WL89);
sram_cell_6t_3 inst_cell_89_81 ( BL81, BLN81, WL89);
sram_cell_6t_3 inst_cell_89_80 ( BL80, BLN80, WL89);
sram_cell_6t_3 inst_cell_89_79 ( BL79, BLN79, WL89);
sram_cell_6t_3 inst_cell_89_78 ( BL78, BLN78, WL89);
sram_cell_6t_3 inst_cell_89_77 ( BL77, BLN77, WL89);
sram_cell_6t_3 inst_cell_89_76 ( BL76, BLN76, WL89);
sram_cell_6t_3 inst_cell_89_75 ( BL75, BLN75, WL89);
sram_cell_6t_3 inst_cell_89_74 ( BL74, BLN74, WL89);
sram_cell_6t_3 inst_cell_89_73 ( BL73, BLN73, WL89);
sram_cell_6t_3 inst_cell_89_72 ( BL72, BLN72, WL89);
sram_cell_6t_3 inst_cell_89_71 ( BL71, BLN71, WL89);
sram_cell_6t_3 inst_cell_89_70 ( BL70, BLN70, WL89);
sram_cell_6t_3 inst_cell_89_69 ( BL69, BLN69, WL89);
sram_cell_6t_3 inst_cell_89_68 ( BL68, BLN68, WL89);
sram_cell_6t_3 inst_cell_89_67 ( BL67, BLN67, WL89);
sram_cell_6t_3 inst_cell_89_66 ( BL66, BLN66, WL89);
sram_cell_6t_3 inst_cell_89_65 ( BL65, BLN65, WL89);
sram_cell_6t_3 inst_cell_89_64 ( BL64, BLN64, WL89);
sram_cell_6t_3 inst_cell_89_63 ( BL63, BLN63, WL89);
sram_cell_6t_3 inst_cell_89_62 ( BL62, BLN62, WL89);
sram_cell_6t_3 inst_cell_89_61 ( BL61, BLN61, WL89);
sram_cell_6t_3 inst_cell_89_60 ( BL60, BLN60, WL89);
sram_cell_6t_3 inst_cell_89_59 ( BL59, BLN59, WL89);
sram_cell_6t_3 inst_cell_89_58 ( BL58, BLN58, WL89);
sram_cell_6t_3 inst_cell_89_57 ( BL57, BLN57, WL89);
sram_cell_6t_3 inst_cell_89_56 ( BL56, BLN56, WL89);
sram_cell_6t_3 inst_cell_89_55 ( BL55, BLN55, WL89);
sram_cell_6t_3 inst_cell_89_54 ( BL54, BLN54, WL89);
sram_cell_6t_3 inst_cell_89_53 ( BL53, BLN53, WL89);
sram_cell_6t_3 inst_cell_89_52 ( BL52, BLN52, WL89);
sram_cell_6t_3 inst_cell_89_51 ( BL51, BLN51, WL89);
sram_cell_6t_3 inst_cell_89_50 ( BL50, BLN50, WL89);
sram_cell_6t_3 inst_cell_89_49 ( BL49, BLN49, WL89);
sram_cell_6t_3 inst_cell_89_48 ( BL48, BLN48, WL89);
sram_cell_6t_3 inst_cell_89_47 ( BL47, BLN47, WL89);
sram_cell_6t_3 inst_cell_89_46 ( BL46, BLN46, WL89);
sram_cell_6t_3 inst_cell_89_45 ( BL45, BLN45, WL89);
sram_cell_6t_3 inst_cell_89_44 ( BL44, BLN44, WL89);
sram_cell_6t_3 inst_cell_89_43 ( BL43, BLN43, WL89);
sram_cell_6t_3 inst_cell_89_42 ( BL42, BLN42, WL89);
sram_cell_6t_3 inst_cell_89_41 ( BL41, BLN41, WL89);
sram_cell_6t_3 inst_cell_89_40 ( BL40, BLN40, WL89);
sram_cell_6t_3 inst_cell_89_39 ( BL39, BLN39, WL89);
sram_cell_6t_3 inst_cell_89_38 ( BL38, BLN38, WL89);
sram_cell_6t_3 inst_cell_89_37 ( BL37, BLN37, WL89);
sram_cell_6t_3 inst_cell_89_36 ( BL36, BLN36, WL89);
sram_cell_6t_3 inst_cell_89_35 ( BL35, BLN35, WL89);
sram_cell_6t_3 inst_cell_89_34 ( BL34, BLN34, WL89);
sram_cell_6t_3 inst_cell_89_33 ( BL33, BLN33, WL89);
sram_cell_6t_3 inst_cell_89_32 ( BL32, BLN32, WL89);
sram_cell_6t_3 inst_cell_89_31 ( BL31, BLN31, WL89);
sram_cell_6t_3 inst_cell_89_30 ( BL30, BLN30, WL89);
sram_cell_6t_3 inst_cell_89_29 ( BL29, BLN29, WL89);
sram_cell_6t_3 inst_cell_89_28 ( BL28, BLN28, WL89);
sram_cell_6t_3 inst_cell_89_27 ( BL27, BLN27, WL89);
sram_cell_6t_3 inst_cell_89_26 ( BL26, BLN26, WL89);
sram_cell_6t_3 inst_cell_89_25 ( BL25, BLN25, WL89);
sram_cell_6t_3 inst_cell_89_24 ( BL24, BLN24, WL89);
sram_cell_6t_3 inst_cell_89_23 ( BL23, BLN23, WL89);
sram_cell_6t_3 inst_cell_89_22 ( BL22, BLN22, WL89);
sram_cell_6t_3 inst_cell_89_21 ( BL21, BLN21, WL89);
sram_cell_6t_3 inst_cell_89_20 ( BL20, BLN20, WL89);
sram_cell_6t_3 inst_cell_89_19 ( BL19, BLN19, WL89);
sram_cell_6t_3 inst_cell_89_18 ( BL18, BLN18, WL89);
sram_cell_6t_3 inst_cell_89_17 ( BL17, BLN17, WL89);
sram_cell_6t_3 inst_cell_89_16 ( BL16, BLN16, WL89);
sram_cell_6t_3 inst_cell_89_15 ( BL15, BLN15, WL89);
sram_cell_6t_3 inst_cell_89_14 ( BL14, BLN14, WL89);
sram_cell_6t_3 inst_cell_89_13 ( BL13, BLN13, WL89);
sram_cell_6t_3 inst_cell_89_12 ( BL12, BLN12, WL89);
sram_cell_6t_3 inst_cell_89_11 ( BL11, BLN11, WL89);
sram_cell_6t_3 inst_cell_89_10 ( BL10, BLN10, WL89);
sram_cell_6t_3 inst_cell_89_9 ( BL9, BLN9, WL89);
sram_cell_6t_3 inst_cell_89_8 ( BL8, BLN8, WL89);
sram_cell_6t_3 inst_cell_89_7 ( BL7, BLN7, WL89);
sram_cell_6t_3 inst_cell_89_6 ( BL6, BLN6, WL89);
sram_cell_6t_3 inst_cell_89_5 ( BL5, BLN5, WL89);
sram_cell_6t_3 inst_cell_89_4 ( BL4, BLN4, WL89);
sram_cell_6t_3 inst_cell_89_3 ( BL3, BLN3, WL89);
sram_cell_6t_3 inst_cell_89_2 ( BL2, BLN2, WL89);
sram_cell_6t_3 inst_cell_89_1 ( BL1, BLN1, WL89);
sram_cell_6t_3 inst_cell_89_0 ( BL0, BLN0, WL89);
sram_cell_6t_3 inst_cell_88_127 ( BL127, BLN127, WL88);
sram_cell_6t_3 inst_cell_88_126 ( BL126, BLN126, WL88);
sram_cell_6t_3 inst_cell_88_125 ( BL125, BLN125, WL88);
sram_cell_6t_3 inst_cell_88_124 ( BL124, BLN124, WL88);
sram_cell_6t_3 inst_cell_88_123 ( BL123, BLN123, WL88);
sram_cell_6t_3 inst_cell_88_122 ( BL122, BLN122, WL88);
sram_cell_6t_3 inst_cell_88_121 ( BL121, BLN121, WL88);
sram_cell_6t_3 inst_cell_88_120 ( BL120, BLN120, WL88);
sram_cell_6t_3 inst_cell_88_119 ( BL119, BLN119, WL88);
sram_cell_6t_3 inst_cell_88_118 ( BL118, BLN118, WL88);
sram_cell_6t_3 inst_cell_88_117 ( BL117, BLN117, WL88);
sram_cell_6t_3 inst_cell_88_116 ( BL116, BLN116, WL88);
sram_cell_6t_3 inst_cell_88_115 ( BL115, BLN115, WL88);
sram_cell_6t_3 inst_cell_88_114 ( BL114, BLN114, WL88);
sram_cell_6t_3 inst_cell_88_113 ( BL113, BLN113, WL88);
sram_cell_6t_3 inst_cell_88_112 ( BL112, BLN112, WL88);
sram_cell_6t_3 inst_cell_88_111 ( BL111, BLN111, WL88);
sram_cell_6t_3 inst_cell_88_110 ( BL110, BLN110, WL88);
sram_cell_6t_3 inst_cell_88_109 ( BL109, BLN109, WL88);
sram_cell_6t_3 inst_cell_88_108 ( BL108, BLN108, WL88);
sram_cell_6t_3 inst_cell_88_107 ( BL107, BLN107, WL88);
sram_cell_6t_3 inst_cell_88_106 ( BL106, BLN106, WL88);
sram_cell_6t_3 inst_cell_88_105 ( BL105, BLN105, WL88);
sram_cell_6t_3 inst_cell_88_104 ( BL104, BLN104, WL88);
sram_cell_6t_3 inst_cell_88_103 ( BL103, BLN103, WL88);
sram_cell_6t_3 inst_cell_88_102 ( BL102, BLN102, WL88);
sram_cell_6t_3 inst_cell_88_101 ( BL101, BLN101, WL88);
sram_cell_6t_3 inst_cell_88_100 ( BL100, BLN100, WL88);
sram_cell_6t_3 inst_cell_88_99 ( BL99, BLN99, WL88);
sram_cell_6t_3 inst_cell_88_98 ( BL98, BLN98, WL88);
sram_cell_6t_3 inst_cell_88_97 ( BL97, BLN97, WL88);
sram_cell_6t_3 inst_cell_88_96 ( BL96, BLN96, WL88);
sram_cell_6t_3 inst_cell_88_95 ( BL95, BLN95, WL88);
sram_cell_6t_3 inst_cell_88_94 ( BL94, BLN94, WL88);
sram_cell_6t_3 inst_cell_88_93 ( BL93, BLN93, WL88);
sram_cell_6t_3 inst_cell_88_92 ( BL92, BLN92, WL88);
sram_cell_6t_3 inst_cell_88_91 ( BL91, BLN91, WL88);
sram_cell_6t_3 inst_cell_88_90 ( BL90, BLN90, WL88);
sram_cell_6t_3 inst_cell_88_89 ( BL89, BLN89, WL88);
sram_cell_6t_3 inst_cell_88_88 ( BL88, BLN88, WL88);
sram_cell_6t_3 inst_cell_88_87 ( BL87, BLN87, WL88);
sram_cell_6t_3 inst_cell_88_86 ( BL86, BLN86, WL88);
sram_cell_6t_3 inst_cell_88_85 ( BL85, BLN85, WL88);
sram_cell_6t_3 inst_cell_88_84 ( BL84, BLN84, WL88);
sram_cell_6t_3 inst_cell_88_83 ( BL83, BLN83, WL88);
sram_cell_6t_3 inst_cell_88_82 ( BL82, BLN82, WL88);
sram_cell_6t_3 inst_cell_88_81 ( BL81, BLN81, WL88);
sram_cell_6t_3 inst_cell_88_80 ( BL80, BLN80, WL88);
sram_cell_6t_3 inst_cell_88_79 ( BL79, BLN79, WL88);
sram_cell_6t_3 inst_cell_88_78 ( BL78, BLN78, WL88);
sram_cell_6t_3 inst_cell_88_77 ( BL77, BLN77, WL88);
sram_cell_6t_3 inst_cell_88_76 ( BL76, BLN76, WL88);
sram_cell_6t_3 inst_cell_88_75 ( BL75, BLN75, WL88);
sram_cell_6t_3 inst_cell_88_74 ( BL74, BLN74, WL88);
sram_cell_6t_3 inst_cell_88_73 ( BL73, BLN73, WL88);
sram_cell_6t_3 inst_cell_88_72 ( BL72, BLN72, WL88);
sram_cell_6t_3 inst_cell_88_71 ( BL71, BLN71, WL88);
sram_cell_6t_3 inst_cell_88_70 ( BL70, BLN70, WL88);
sram_cell_6t_3 inst_cell_88_69 ( BL69, BLN69, WL88);
sram_cell_6t_3 inst_cell_88_68 ( BL68, BLN68, WL88);
sram_cell_6t_3 inst_cell_88_67 ( BL67, BLN67, WL88);
sram_cell_6t_3 inst_cell_88_66 ( BL66, BLN66, WL88);
sram_cell_6t_3 inst_cell_88_65 ( BL65, BLN65, WL88);
sram_cell_6t_3 inst_cell_88_64 ( BL64, BLN64, WL88);
sram_cell_6t_3 inst_cell_88_63 ( BL63, BLN63, WL88);
sram_cell_6t_3 inst_cell_88_62 ( BL62, BLN62, WL88);
sram_cell_6t_3 inst_cell_88_61 ( BL61, BLN61, WL88);
sram_cell_6t_3 inst_cell_88_60 ( BL60, BLN60, WL88);
sram_cell_6t_3 inst_cell_88_59 ( BL59, BLN59, WL88);
sram_cell_6t_3 inst_cell_88_58 ( BL58, BLN58, WL88);
sram_cell_6t_3 inst_cell_88_57 ( BL57, BLN57, WL88);
sram_cell_6t_3 inst_cell_88_56 ( BL56, BLN56, WL88);
sram_cell_6t_3 inst_cell_88_55 ( BL55, BLN55, WL88);
sram_cell_6t_3 inst_cell_88_54 ( BL54, BLN54, WL88);
sram_cell_6t_3 inst_cell_88_53 ( BL53, BLN53, WL88);
sram_cell_6t_3 inst_cell_88_52 ( BL52, BLN52, WL88);
sram_cell_6t_3 inst_cell_88_51 ( BL51, BLN51, WL88);
sram_cell_6t_3 inst_cell_88_50 ( BL50, BLN50, WL88);
sram_cell_6t_3 inst_cell_88_49 ( BL49, BLN49, WL88);
sram_cell_6t_3 inst_cell_88_48 ( BL48, BLN48, WL88);
sram_cell_6t_3 inst_cell_88_47 ( BL47, BLN47, WL88);
sram_cell_6t_3 inst_cell_88_46 ( BL46, BLN46, WL88);
sram_cell_6t_3 inst_cell_88_45 ( BL45, BLN45, WL88);
sram_cell_6t_3 inst_cell_88_44 ( BL44, BLN44, WL88);
sram_cell_6t_3 inst_cell_88_43 ( BL43, BLN43, WL88);
sram_cell_6t_3 inst_cell_88_42 ( BL42, BLN42, WL88);
sram_cell_6t_3 inst_cell_88_41 ( BL41, BLN41, WL88);
sram_cell_6t_3 inst_cell_88_40 ( BL40, BLN40, WL88);
sram_cell_6t_3 inst_cell_88_39 ( BL39, BLN39, WL88);
sram_cell_6t_3 inst_cell_88_38 ( BL38, BLN38, WL88);
sram_cell_6t_3 inst_cell_88_37 ( BL37, BLN37, WL88);
sram_cell_6t_3 inst_cell_88_36 ( BL36, BLN36, WL88);
sram_cell_6t_3 inst_cell_88_35 ( BL35, BLN35, WL88);
sram_cell_6t_3 inst_cell_88_34 ( BL34, BLN34, WL88);
sram_cell_6t_3 inst_cell_88_33 ( BL33, BLN33, WL88);
sram_cell_6t_3 inst_cell_88_32 ( BL32, BLN32, WL88);
sram_cell_6t_3 inst_cell_88_31 ( BL31, BLN31, WL88);
sram_cell_6t_3 inst_cell_88_30 ( BL30, BLN30, WL88);
sram_cell_6t_3 inst_cell_88_29 ( BL29, BLN29, WL88);
sram_cell_6t_3 inst_cell_88_28 ( BL28, BLN28, WL88);
sram_cell_6t_3 inst_cell_88_27 ( BL27, BLN27, WL88);
sram_cell_6t_3 inst_cell_88_26 ( BL26, BLN26, WL88);
sram_cell_6t_3 inst_cell_88_25 ( BL25, BLN25, WL88);
sram_cell_6t_3 inst_cell_88_24 ( BL24, BLN24, WL88);
sram_cell_6t_3 inst_cell_88_23 ( BL23, BLN23, WL88);
sram_cell_6t_3 inst_cell_88_22 ( BL22, BLN22, WL88);
sram_cell_6t_3 inst_cell_88_21 ( BL21, BLN21, WL88);
sram_cell_6t_3 inst_cell_88_20 ( BL20, BLN20, WL88);
sram_cell_6t_3 inst_cell_88_19 ( BL19, BLN19, WL88);
sram_cell_6t_3 inst_cell_88_18 ( BL18, BLN18, WL88);
sram_cell_6t_3 inst_cell_88_17 ( BL17, BLN17, WL88);
sram_cell_6t_3 inst_cell_88_16 ( BL16, BLN16, WL88);
sram_cell_6t_3 inst_cell_88_15 ( BL15, BLN15, WL88);
sram_cell_6t_3 inst_cell_88_14 ( BL14, BLN14, WL88);
sram_cell_6t_3 inst_cell_88_13 ( BL13, BLN13, WL88);
sram_cell_6t_3 inst_cell_88_12 ( BL12, BLN12, WL88);
sram_cell_6t_3 inst_cell_88_11 ( BL11, BLN11, WL88);
sram_cell_6t_3 inst_cell_88_10 ( BL10, BLN10, WL88);
sram_cell_6t_3 inst_cell_88_9 ( BL9, BLN9, WL88);
sram_cell_6t_3 inst_cell_88_8 ( BL8, BLN8, WL88);
sram_cell_6t_3 inst_cell_88_7 ( BL7, BLN7, WL88);
sram_cell_6t_3 inst_cell_88_6 ( BL6, BLN6, WL88);
sram_cell_6t_3 inst_cell_88_5 ( BL5, BLN5, WL88);
sram_cell_6t_3 inst_cell_88_4 ( BL4, BLN4, WL88);
sram_cell_6t_3 inst_cell_88_3 ( BL3, BLN3, WL88);
sram_cell_6t_3 inst_cell_88_2 ( BL2, BLN2, WL88);
sram_cell_6t_3 inst_cell_88_1 ( BL1, BLN1, WL88);
sram_cell_6t_3 inst_cell_88_0 ( BL0, BLN0, WL88);
sram_cell_6t_3 inst_cell_87_127 ( BL127, BLN127, WL87);
sram_cell_6t_3 inst_cell_87_126 ( BL126, BLN126, WL87);
sram_cell_6t_3 inst_cell_87_125 ( BL125, BLN125, WL87);
sram_cell_6t_3 inst_cell_87_124 ( BL124, BLN124, WL87);
sram_cell_6t_3 inst_cell_87_123 ( BL123, BLN123, WL87);
sram_cell_6t_3 inst_cell_87_122 ( BL122, BLN122, WL87);
sram_cell_6t_3 inst_cell_87_121 ( BL121, BLN121, WL87);
sram_cell_6t_3 inst_cell_87_120 ( BL120, BLN120, WL87);
sram_cell_6t_3 inst_cell_87_119 ( BL119, BLN119, WL87);
sram_cell_6t_3 inst_cell_87_118 ( BL118, BLN118, WL87);
sram_cell_6t_3 inst_cell_87_117 ( BL117, BLN117, WL87);
sram_cell_6t_3 inst_cell_87_116 ( BL116, BLN116, WL87);
sram_cell_6t_3 inst_cell_87_115 ( BL115, BLN115, WL87);
sram_cell_6t_3 inst_cell_87_114 ( BL114, BLN114, WL87);
sram_cell_6t_3 inst_cell_87_113 ( BL113, BLN113, WL87);
sram_cell_6t_3 inst_cell_87_112 ( BL112, BLN112, WL87);
sram_cell_6t_3 inst_cell_87_111 ( BL111, BLN111, WL87);
sram_cell_6t_3 inst_cell_87_110 ( BL110, BLN110, WL87);
sram_cell_6t_3 inst_cell_87_109 ( BL109, BLN109, WL87);
sram_cell_6t_3 inst_cell_87_108 ( BL108, BLN108, WL87);
sram_cell_6t_3 inst_cell_87_107 ( BL107, BLN107, WL87);
sram_cell_6t_3 inst_cell_87_106 ( BL106, BLN106, WL87);
sram_cell_6t_3 inst_cell_87_105 ( BL105, BLN105, WL87);
sram_cell_6t_3 inst_cell_87_104 ( BL104, BLN104, WL87);
sram_cell_6t_3 inst_cell_87_103 ( BL103, BLN103, WL87);
sram_cell_6t_3 inst_cell_87_102 ( BL102, BLN102, WL87);
sram_cell_6t_3 inst_cell_87_101 ( BL101, BLN101, WL87);
sram_cell_6t_3 inst_cell_87_100 ( BL100, BLN100, WL87);
sram_cell_6t_3 inst_cell_87_99 ( BL99, BLN99, WL87);
sram_cell_6t_3 inst_cell_87_98 ( BL98, BLN98, WL87);
sram_cell_6t_3 inst_cell_87_97 ( BL97, BLN97, WL87);
sram_cell_6t_3 inst_cell_87_96 ( BL96, BLN96, WL87);
sram_cell_6t_3 inst_cell_87_95 ( BL95, BLN95, WL87);
sram_cell_6t_3 inst_cell_87_94 ( BL94, BLN94, WL87);
sram_cell_6t_3 inst_cell_87_93 ( BL93, BLN93, WL87);
sram_cell_6t_3 inst_cell_87_92 ( BL92, BLN92, WL87);
sram_cell_6t_3 inst_cell_87_91 ( BL91, BLN91, WL87);
sram_cell_6t_3 inst_cell_87_90 ( BL90, BLN90, WL87);
sram_cell_6t_3 inst_cell_87_89 ( BL89, BLN89, WL87);
sram_cell_6t_3 inst_cell_87_88 ( BL88, BLN88, WL87);
sram_cell_6t_3 inst_cell_87_87 ( BL87, BLN87, WL87);
sram_cell_6t_3 inst_cell_87_86 ( BL86, BLN86, WL87);
sram_cell_6t_3 inst_cell_87_85 ( BL85, BLN85, WL87);
sram_cell_6t_3 inst_cell_87_84 ( BL84, BLN84, WL87);
sram_cell_6t_3 inst_cell_87_83 ( BL83, BLN83, WL87);
sram_cell_6t_3 inst_cell_87_82 ( BL82, BLN82, WL87);
sram_cell_6t_3 inst_cell_87_81 ( BL81, BLN81, WL87);
sram_cell_6t_3 inst_cell_87_80 ( BL80, BLN80, WL87);
sram_cell_6t_3 inst_cell_87_79 ( BL79, BLN79, WL87);
sram_cell_6t_3 inst_cell_87_78 ( BL78, BLN78, WL87);
sram_cell_6t_3 inst_cell_87_77 ( BL77, BLN77, WL87);
sram_cell_6t_3 inst_cell_87_76 ( BL76, BLN76, WL87);
sram_cell_6t_3 inst_cell_87_75 ( BL75, BLN75, WL87);
sram_cell_6t_3 inst_cell_87_74 ( BL74, BLN74, WL87);
sram_cell_6t_3 inst_cell_87_73 ( BL73, BLN73, WL87);
sram_cell_6t_3 inst_cell_87_72 ( BL72, BLN72, WL87);
sram_cell_6t_3 inst_cell_87_71 ( BL71, BLN71, WL87);
sram_cell_6t_3 inst_cell_87_70 ( BL70, BLN70, WL87);
sram_cell_6t_3 inst_cell_87_69 ( BL69, BLN69, WL87);
sram_cell_6t_3 inst_cell_87_68 ( BL68, BLN68, WL87);
sram_cell_6t_3 inst_cell_87_67 ( BL67, BLN67, WL87);
sram_cell_6t_3 inst_cell_87_66 ( BL66, BLN66, WL87);
sram_cell_6t_3 inst_cell_87_65 ( BL65, BLN65, WL87);
sram_cell_6t_3 inst_cell_87_64 ( BL64, BLN64, WL87);
sram_cell_6t_3 inst_cell_87_63 ( BL63, BLN63, WL87);
sram_cell_6t_3 inst_cell_87_62 ( BL62, BLN62, WL87);
sram_cell_6t_3 inst_cell_87_61 ( BL61, BLN61, WL87);
sram_cell_6t_3 inst_cell_87_60 ( BL60, BLN60, WL87);
sram_cell_6t_3 inst_cell_87_59 ( BL59, BLN59, WL87);
sram_cell_6t_3 inst_cell_87_58 ( BL58, BLN58, WL87);
sram_cell_6t_3 inst_cell_87_57 ( BL57, BLN57, WL87);
sram_cell_6t_3 inst_cell_87_56 ( BL56, BLN56, WL87);
sram_cell_6t_3 inst_cell_87_55 ( BL55, BLN55, WL87);
sram_cell_6t_3 inst_cell_87_54 ( BL54, BLN54, WL87);
sram_cell_6t_3 inst_cell_87_53 ( BL53, BLN53, WL87);
sram_cell_6t_3 inst_cell_87_52 ( BL52, BLN52, WL87);
sram_cell_6t_3 inst_cell_87_51 ( BL51, BLN51, WL87);
sram_cell_6t_3 inst_cell_87_50 ( BL50, BLN50, WL87);
sram_cell_6t_3 inst_cell_87_49 ( BL49, BLN49, WL87);
sram_cell_6t_3 inst_cell_87_48 ( BL48, BLN48, WL87);
sram_cell_6t_3 inst_cell_87_47 ( BL47, BLN47, WL87);
sram_cell_6t_3 inst_cell_87_46 ( BL46, BLN46, WL87);
sram_cell_6t_3 inst_cell_87_45 ( BL45, BLN45, WL87);
sram_cell_6t_3 inst_cell_87_44 ( BL44, BLN44, WL87);
sram_cell_6t_3 inst_cell_87_43 ( BL43, BLN43, WL87);
sram_cell_6t_3 inst_cell_87_42 ( BL42, BLN42, WL87);
sram_cell_6t_3 inst_cell_87_41 ( BL41, BLN41, WL87);
sram_cell_6t_3 inst_cell_87_40 ( BL40, BLN40, WL87);
sram_cell_6t_3 inst_cell_87_39 ( BL39, BLN39, WL87);
sram_cell_6t_3 inst_cell_87_38 ( BL38, BLN38, WL87);
sram_cell_6t_3 inst_cell_87_37 ( BL37, BLN37, WL87);
sram_cell_6t_3 inst_cell_87_36 ( BL36, BLN36, WL87);
sram_cell_6t_3 inst_cell_87_35 ( BL35, BLN35, WL87);
sram_cell_6t_3 inst_cell_87_34 ( BL34, BLN34, WL87);
sram_cell_6t_3 inst_cell_87_33 ( BL33, BLN33, WL87);
sram_cell_6t_3 inst_cell_87_32 ( BL32, BLN32, WL87);
sram_cell_6t_3 inst_cell_87_31 ( BL31, BLN31, WL87);
sram_cell_6t_3 inst_cell_87_30 ( BL30, BLN30, WL87);
sram_cell_6t_3 inst_cell_87_29 ( BL29, BLN29, WL87);
sram_cell_6t_3 inst_cell_87_28 ( BL28, BLN28, WL87);
sram_cell_6t_3 inst_cell_87_27 ( BL27, BLN27, WL87);
sram_cell_6t_3 inst_cell_87_26 ( BL26, BLN26, WL87);
sram_cell_6t_3 inst_cell_87_25 ( BL25, BLN25, WL87);
sram_cell_6t_3 inst_cell_87_24 ( BL24, BLN24, WL87);
sram_cell_6t_3 inst_cell_87_23 ( BL23, BLN23, WL87);
sram_cell_6t_3 inst_cell_87_22 ( BL22, BLN22, WL87);
sram_cell_6t_3 inst_cell_87_21 ( BL21, BLN21, WL87);
sram_cell_6t_3 inst_cell_87_20 ( BL20, BLN20, WL87);
sram_cell_6t_3 inst_cell_87_19 ( BL19, BLN19, WL87);
sram_cell_6t_3 inst_cell_87_18 ( BL18, BLN18, WL87);
sram_cell_6t_3 inst_cell_87_17 ( BL17, BLN17, WL87);
sram_cell_6t_3 inst_cell_87_16 ( BL16, BLN16, WL87);
sram_cell_6t_3 inst_cell_87_15 ( BL15, BLN15, WL87);
sram_cell_6t_3 inst_cell_87_14 ( BL14, BLN14, WL87);
sram_cell_6t_3 inst_cell_87_13 ( BL13, BLN13, WL87);
sram_cell_6t_3 inst_cell_87_12 ( BL12, BLN12, WL87);
sram_cell_6t_3 inst_cell_87_11 ( BL11, BLN11, WL87);
sram_cell_6t_3 inst_cell_87_10 ( BL10, BLN10, WL87);
sram_cell_6t_3 inst_cell_87_9 ( BL9, BLN9, WL87);
sram_cell_6t_3 inst_cell_87_8 ( BL8, BLN8, WL87);
sram_cell_6t_3 inst_cell_87_7 ( BL7, BLN7, WL87);
sram_cell_6t_3 inst_cell_87_6 ( BL6, BLN6, WL87);
sram_cell_6t_3 inst_cell_87_5 ( BL5, BLN5, WL87);
sram_cell_6t_3 inst_cell_87_4 ( BL4, BLN4, WL87);
sram_cell_6t_3 inst_cell_87_3 ( BL3, BLN3, WL87);
sram_cell_6t_3 inst_cell_87_2 ( BL2, BLN2, WL87);
sram_cell_6t_3 inst_cell_87_1 ( BL1, BLN1, WL87);
sram_cell_6t_3 inst_cell_87_0 ( BL0, BLN0, WL87);
sram_cell_6t_3 inst_cell_86_127 ( BL127, BLN127, WL86);
sram_cell_6t_3 inst_cell_86_126 ( BL126, BLN126, WL86);
sram_cell_6t_3 inst_cell_86_125 ( BL125, BLN125, WL86);
sram_cell_6t_3 inst_cell_86_124 ( BL124, BLN124, WL86);
sram_cell_6t_3 inst_cell_86_123 ( BL123, BLN123, WL86);
sram_cell_6t_3 inst_cell_86_122 ( BL122, BLN122, WL86);
sram_cell_6t_3 inst_cell_86_121 ( BL121, BLN121, WL86);
sram_cell_6t_3 inst_cell_86_120 ( BL120, BLN120, WL86);
sram_cell_6t_3 inst_cell_86_119 ( BL119, BLN119, WL86);
sram_cell_6t_3 inst_cell_86_118 ( BL118, BLN118, WL86);
sram_cell_6t_3 inst_cell_86_117 ( BL117, BLN117, WL86);
sram_cell_6t_3 inst_cell_86_116 ( BL116, BLN116, WL86);
sram_cell_6t_3 inst_cell_86_115 ( BL115, BLN115, WL86);
sram_cell_6t_3 inst_cell_86_114 ( BL114, BLN114, WL86);
sram_cell_6t_3 inst_cell_86_113 ( BL113, BLN113, WL86);
sram_cell_6t_3 inst_cell_86_112 ( BL112, BLN112, WL86);
sram_cell_6t_3 inst_cell_86_111 ( BL111, BLN111, WL86);
sram_cell_6t_3 inst_cell_86_110 ( BL110, BLN110, WL86);
sram_cell_6t_3 inst_cell_86_109 ( BL109, BLN109, WL86);
sram_cell_6t_3 inst_cell_86_108 ( BL108, BLN108, WL86);
sram_cell_6t_3 inst_cell_86_107 ( BL107, BLN107, WL86);
sram_cell_6t_3 inst_cell_86_106 ( BL106, BLN106, WL86);
sram_cell_6t_3 inst_cell_86_105 ( BL105, BLN105, WL86);
sram_cell_6t_3 inst_cell_86_104 ( BL104, BLN104, WL86);
sram_cell_6t_3 inst_cell_86_103 ( BL103, BLN103, WL86);
sram_cell_6t_3 inst_cell_86_102 ( BL102, BLN102, WL86);
sram_cell_6t_3 inst_cell_86_101 ( BL101, BLN101, WL86);
sram_cell_6t_3 inst_cell_86_100 ( BL100, BLN100, WL86);
sram_cell_6t_3 inst_cell_86_99 ( BL99, BLN99, WL86);
sram_cell_6t_3 inst_cell_86_98 ( BL98, BLN98, WL86);
sram_cell_6t_3 inst_cell_86_97 ( BL97, BLN97, WL86);
sram_cell_6t_3 inst_cell_86_96 ( BL96, BLN96, WL86);
sram_cell_6t_3 inst_cell_86_95 ( BL95, BLN95, WL86);
sram_cell_6t_3 inst_cell_86_94 ( BL94, BLN94, WL86);
sram_cell_6t_3 inst_cell_86_93 ( BL93, BLN93, WL86);
sram_cell_6t_3 inst_cell_86_92 ( BL92, BLN92, WL86);
sram_cell_6t_3 inst_cell_86_91 ( BL91, BLN91, WL86);
sram_cell_6t_3 inst_cell_86_90 ( BL90, BLN90, WL86);
sram_cell_6t_3 inst_cell_86_89 ( BL89, BLN89, WL86);
sram_cell_6t_3 inst_cell_86_88 ( BL88, BLN88, WL86);
sram_cell_6t_3 inst_cell_86_87 ( BL87, BLN87, WL86);
sram_cell_6t_3 inst_cell_86_86 ( BL86, BLN86, WL86);
sram_cell_6t_3 inst_cell_86_85 ( BL85, BLN85, WL86);
sram_cell_6t_3 inst_cell_86_84 ( BL84, BLN84, WL86);
sram_cell_6t_3 inst_cell_86_83 ( BL83, BLN83, WL86);
sram_cell_6t_3 inst_cell_86_82 ( BL82, BLN82, WL86);
sram_cell_6t_3 inst_cell_86_81 ( BL81, BLN81, WL86);
sram_cell_6t_3 inst_cell_86_80 ( BL80, BLN80, WL86);
sram_cell_6t_3 inst_cell_86_79 ( BL79, BLN79, WL86);
sram_cell_6t_3 inst_cell_86_78 ( BL78, BLN78, WL86);
sram_cell_6t_3 inst_cell_86_77 ( BL77, BLN77, WL86);
sram_cell_6t_3 inst_cell_86_76 ( BL76, BLN76, WL86);
sram_cell_6t_3 inst_cell_86_75 ( BL75, BLN75, WL86);
sram_cell_6t_3 inst_cell_86_74 ( BL74, BLN74, WL86);
sram_cell_6t_3 inst_cell_86_73 ( BL73, BLN73, WL86);
sram_cell_6t_3 inst_cell_86_72 ( BL72, BLN72, WL86);
sram_cell_6t_3 inst_cell_86_71 ( BL71, BLN71, WL86);
sram_cell_6t_3 inst_cell_86_70 ( BL70, BLN70, WL86);
sram_cell_6t_3 inst_cell_86_69 ( BL69, BLN69, WL86);
sram_cell_6t_3 inst_cell_86_68 ( BL68, BLN68, WL86);
sram_cell_6t_3 inst_cell_86_67 ( BL67, BLN67, WL86);
sram_cell_6t_3 inst_cell_86_66 ( BL66, BLN66, WL86);
sram_cell_6t_3 inst_cell_86_65 ( BL65, BLN65, WL86);
sram_cell_6t_3 inst_cell_86_64 ( BL64, BLN64, WL86);
sram_cell_6t_3 inst_cell_86_63 ( BL63, BLN63, WL86);
sram_cell_6t_3 inst_cell_86_62 ( BL62, BLN62, WL86);
sram_cell_6t_3 inst_cell_86_61 ( BL61, BLN61, WL86);
sram_cell_6t_3 inst_cell_86_60 ( BL60, BLN60, WL86);
sram_cell_6t_3 inst_cell_86_59 ( BL59, BLN59, WL86);
sram_cell_6t_3 inst_cell_86_58 ( BL58, BLN58, WL86);
sram_cell_6t_3 inst_cell_86_57 ( BL57, BLN57, WL86);
sram_cell_6t_3 inst_cell_86_56 ( BL56, BLN56, WL86);
sram_cell_6t_3 inst_cell_86_55 ( BL55, BLN55, WL86);
sram_cell_6t_3 inst_cell_86_54 ( BL54, BLN54, WL86);
sram_cell_6t_3 inst_cell_86_53 ( BL53, BLN53, WL86);
sram_cell_6t_3 inst_cell_86_52 ( BL52, BLN52, WL86);
sram_cell_6t_3 inst_cell_86_51 ( BL51, BLN51, WL86);
sram_cell_6t_3 inst_cell_86_50 ( BL50, BLN50, WL86);
sram_cell_6t_3 inst_cell_86_49 ( BL49, BLN49, WL86);
sram_cell_6t_3 inst_cell_86_48 ( BL48, BLN48, WL86);
sram_cell_6t_3 inst_cell_86_47 ( BL47, BLN47, WL86);
sram_cell_6t_3 inst_cell_86_46 ( BL46, BLN46, WL86);
sram_cell_6t_3 inst_cell_86_45 ( BL45, BLN45, WL86);
sram_cell_6t_3 inst_cell_86_44 ( BL44, BLN44, WL86);
sram_cell_6t_3 inst_cell_86_43 ( BL43, BLN43, WL86);
sram_cell_6t_3 inst_cell_86_42 ( BL42, BLN42, WL86);
sram_cell_6t_3 inst_cell_86_41 ( BL41, BLN41, WL86);
sram_cell_6t_3 inst_cell_86_40 ( BL40, BLN40, WL86);
sram_cell_6t_3 inst_cell_86_39 ( BL39, BLN39, WL86);
sram_cell_6t_3 inst_cell_86_38 ( BL38, BLN38, WL86);
sram_cell_6t_3 inst_cell_86_37 ( BL37, BLN37, WL86);
sram_cell_6t_3 inst_cell_86_36 ( BL36, BLN36, WL86);
sram_cell_6t_3 inst_cell_86_35 ( BL35, BLN35, WL86);
sram_cell_6t_3 inst_cell_86_34 ( BL34, BLN34, WL86);
sram_cell_6t_3 inst_cell_86_33 ( BL33, BLN33, WL86);
sram_cell_6t_3 inst_cell_86_32 ( BL32, BLN32, WL86);
sram_cell_6t_3 inst_cell_86_31 ( BL31, BLN31, WL86);
sram_cell_6t_3 inst_cell_86_30 ( BL30, BLN30, WL86);
sram_cell_6t_3 inst_cell_86_29 ( BL29, BLN29, WL86);
sram_cell_6t_3 inst_cell_86_28 ( BL28, BLN28, WL86);
sram_cell_6t_3 inst_cell_86_27 ( BL27, BLN27, WL86);
sram_cell_6t_3 inst_cell_86_26 ( BL26, BLN26, WL86);
sram_cell_6t_3 inst_cell_86_25 ( BL25, BLN25, WL86);
sram_cell_6t_3 inst_cell_86_24 ( BL24, BLN24, WL86);
sram_cell_6t_3 inst_cell_86_23 ( BL23, BLN23, WL86);
sram_cell_6t_3 inst_cell_86_22 ( BL22, BLN22, WL86);
sram_cell_6t_3 inst_cell_86_21 ( BL21, BLN21, WL86);
sram_cell_6t_3 inst_cell_86_20 ( BL20, BLN20, WL86);
sram_cell_6t_3 inst_cell_86_19 ( BL19, BLN19, WL86);
sram_cell_6t_3 inst_cell_86_18 ( BL18, BLN18, WL86);
sram_cell_6t_3 inst_cell_86_17 ( BL17, BLN17, WL86);
sram_cell_6t_3 inst_cell_86_16 ( BL16, BLN16, WL86);
sram_cell_6t_3 inst_cell_86_15 ( BL15, BLN15, WL86);
sram_cell_6t_3 inst_cell_86_14 ( BL14, BLN14, WL86);
sram_cell_6t_3 inst_cell_86_13 ( BL13, BLN13, WL86);
sram_cell_6t_3 inst_cell_86_12 ( BL12, BLN12, WL86);
sram_cell_6t_3 inst_cell_86_11 ( BL11, BLN11, WL86);
sram_cell_6t_3 inst_cell_86_10 ( BL10, BLN10, WL86);
sram_cell_6t_3 inst_cell_86_9 ( BL9, BLN9, WL86);
sram_cell_6t_3 inst_cell_86_8 ( BL8, BLN8, WL86);
sram_cell_6t_3 inst_cell_86_7 ( BL7, BLN7, WL86);
sram_cell_6t_3 inst_cell_86_6 ( BL6, BLN6, WL86);
sram_cell_6t_3 inst_cell_86_5 ( BL5, BLN5, WL86);
sram_cell_6t_3 inst_cell_86_4 ( BL4, BLN4, WL86);
sram_cell_6t_3 inst_cell_86_3 ( BL3, BLN3, WL86);
sram_cell_6t_3 inst_cell_86_2 ( BL2, BLN2, WL86);
sram_cell_6t_3 inst_cell_86_1 ( BL1, BLN1, WL86);
sram_cell_6t_3 inst_cell_86_0 ( BL0, BLN0, WL86);
sram_cell_6t_3 inst_cell_85_127 ( BL127, BLN127, WL85);
sram_cell_6t_3 inst_cell_85_126 ( BL126, BLN126, WL85);
sram_cell_6t_3 inst_cell_85_125 ( BL125, BLN125, WL85);
sram_cell_6t_3 inst_cell_85_124 ( BL124, BLN124, WL85);
sram_cell_6t_3 inst_cell_85_123 ( BL123, BLN123, WL85);
sram_cell_6t_3 inst_cell_85_122 ( BL122, BLN122, WL85);
sram_cell_6t_3 inst_cell_85_121 ( BL121, BLN121, WL85);
sram_cell_6t_3 inst_cell_85_120 ( BL120, BLN120, WL85);
sram_cell_6t_3 inst_cell_85_119 ( BL119, BLN119, WL85);
sram_cell_6t_3 inst_cell_85_118 ( BL118, BLN118, WL85);
sram_cell_6t_3 inst_cell_85_117 ( BL117, BLN117, WL85);
sram_cell_6t_3 inst_cell_85_116 ( BL116, BLN116, WL85);
sram_cell_6t_3 inst_cell_85_115 ( BL115, BLN115, WL85);
sram_cell_6t_3 inst_cell_85_114 ( BL114, BLN114, WL85);
sram_cell_6t_3 inst_cell_85_113 ( BL113, BLN113, WL85);
sram_cell_6t_3 inst_cell_85_112 ( BL112, BLN112, WL85);
sram_cell_6t_3 inst_cell_85_111 ( BL111, BLN111, WL85);
sram_cell_6t_3 inst_cell_85_110 ( BL110, BLN110, WL85);
sram_cell_6t_3 inst_cell_85_109 ( BL109, BLN109, WL85);
sram_cell_6t_3 inst_cell_85_108 ( BL108, BLN108, WL85);
sram_cell_6t_3 inst_cell_85_107 ( BL107, BLN107, WL85);
sram_cell_6t_3 inst_cell_85_106 ( BL106, BLN106, WL85);
sram_cell_6t_3 inst_cell_85_105 ( BL105, BLN105, WL85);
sram_cell_6t_3 inst_cell_85_104 ( BL104, BLN104, WL85);
sram_cell_6t_3 inst_cell_85_103 ( BL103, BLN103, WL85);
sram_cell_6t_3 inst_cell_85_102 ( BL102, BLN102, WL85);
sram_cell_6t_3 inst_cell_85_101 ( BL101, BLN101, WL85);
sram_cell_6t_3 inst_cell_85_100 ( BL100, BLN100, WL85);
sram_cell_6t_3 inst_cell_85_99 ( BL99, BLN99, WL85);
sram_cell_6t_3 inst_cell_85_98 ( BL98, BLN98, WL85);
sram_cell_6t_3 inst_cell_85_97 ( BL97, BLN97, WL85);
sram_cell_6t_3 inst_cell_85_96 ( BL96, BLN96, WL85);
sram_cell_6t_3 inst_cell_85_95 ( BL95, BLN95, WL85);
sram_cell_6t_3 inst_cell_85_94 ( BL94, BLN94, WL85);
sram_cell_6t_3 inst_cell_85_93 ( BL93, BLN93, WL85);
sram_cell_6t_3 inst_cell_85_92 ( BL92, BLN92, WL85);
sram_cell_6t_3 inst_cell_85_91 ( BL91, BLN91, WL85);
sram_cell_6t_3 inst_cell_85_90 ( BL90, BLN90, WL85);
sram_cell_6t_3 inst_cell_85_89 ( BL89, BLN89, WL85);
sram_cell_6t_3 inst_cell_85_88 ( BL88, BLN88, WL85);
sram_cell_6t_3 inst_cell_85_87 ( BL87, BLN87, WL85);
sram_cell_6t_3 inst_cell_85_86 ( BL86, BLN86, WL85);
sram_cell_6t_3 inst_cell_85_85 ( BL85, BLN85, WL85);
sram_cell_6t_3 inst_cell_85_84 ( BL84, BLN84, WL85);
sram_cell_6t_3 inst_cell_85_83 ( BL83, BLN83, WL85);
sram_cell_6t_3 inst_cell_85_82 ( BL82, BLN82, WL85);
sram_cell_6t_3 inst_cell_85_81 ( BL81, BLN81, WL85);
sram_cell_6t_3 inst_cell_85_80 ( BL80, BLN80, WL85);
sram_cell_6t_3 inst_cell_85_79 ( BL79, BLN79, WL85);
sram_cell_6t_3 inst_cell_85_78 ( BL78, BLN78, WL85);
sram_cell_6t_3 inst_cell_85_77 ( BL77, BLN77, WL85);
sram_cell_6t_3 inst_cell_85_76 ( BL76, BLN76, WL85);
sram_cell_6t_3 inst_cell_85_75 ( BL75, BLN75, WL85);
sram_cell_6t_3 inst_cell_85_74 ( BL74, BLN74, WL85);
sram_cell_6t_3 inst_cell_85_73 ( BL73, BLN73, WL85);
sram_cell_6t_3 inst_cell_85_72 ( BL72, BLN72, WL85);
sram_cell_6t_3 inst_cell_85_71 ( BL71, BLN71, WL85);
sram_cell_6t_3 inst_cell_85_70 ( BL70, BLN70, WL85);
sram_cell_6t_3 inst_cell_85_69 ( BL69, BLN69, WL85);
sram_cell_6t_3 inst_cell_85_68 ( BL68, BLN68, WL85);
sram_cell_6t_3 inst_cell_85_67 ( BL67, BLN67, WL85);
sram_cell_6t_3 inst_cell_85_66 ( BL66, BLN66, WL85);
sram_cell_6t_3 inst_cell_85_65 ( BL65, BLN65, WL85);
sram_cell_6t_3 inst_cell_85_64 ( BL64, BLN64, WL85);
sram_cell_6t_3 inst_cell_85_63 ( BL63, BLN63, WL85);
sram_cell_6t_3 inst_cell_85_62 ( BL62, BLN62, WL85);
sram_cell_6t_3 inst_cell_85_61 ( BL61, BLN61, WL85);
sram_cell_6t_3 inst_cell_85_60 ( BL60, BLN60, WL85);
sram_cell_6t_3 inst_cell_85_59 ( BL59, BLN59, WL85);
sram_cell_6t_3 inst_cell_85_58 ( BL58, BLN58, WL85);
sram_cell_6t_3 inst_cell_85_57 ( BL57, BLN57, WL85);
sram_cell_6t_3 inst_cell_85_56 ( BL56, BLN56, WL85);
sram_cell_6t_3 inst_cell_85_55 ( BL55, BLN55, WL85);
sram_cell_6t_3 inst_cell_85_54 ( BL54, BLN54, WL85);
sram_cell_6t_3 inst_cell_85_53 ( BL53, BLN53, WL85);
sram_cell_6t_3 inst_cell_85_52 ( BL52, BLN52, WL85);
sram_cell_6t_3 inst_cell_85_51 ( BL51, BLN51, WL85);
sram_cell_6t_3 inst_cell_85_50 ( BL50, BLN50, WL85);
sram_cell_6t_3 inst_cell_85_49 ( BL49, BLN49, WL85);
sram_cell_6t_3 inst_cell_85_48 ( BL48, BLN48, WL85);
sram_cell_6t_3 inst_cell_85_47 ( BL47, BLN47, WL85);
sram_cell_6t_3 inst_cell_85_46 ( BL46, BLN46, WL85);
sram_cell_6t_3 inst_cell_85_45 ( BL45, BLN45, WL85);
sram_cell_6t_3 inst_cell_85_44 ( BL44, BLN44, WL85);
sram_cell_6t_3 inst_cell_85_43 ( BL43, BLN43, WL85);
sram_cell_6t_3 inst_cell_85_42 ( BL42, BLN42, WL85);
sram_cell_6t_3 inst_cell_85_41 ( BL41, BLN41, WL85);
sram_cell_6t_3 inst_cell_85_40 ( BL40, BLN40, WL85);
sram_cell_6t_3 inst_cell_85_39 ( BL39, BLN39, WL85);
sram_cell_6t_3 inst_cell_85_38 ( BL38, BLN38, WL85);
sram_cell_6t_3 inst_cell_85_37 ( BL37, BLN37, WL85);
sram_cell_6t_3 inst_cell_85_36 ( BL36, BLN36, WL85);
sram_cell_6t_3 inst_cell_85_35 ( BL35, BLN35, WL85);
sram_cell_6t_3 inst_cell_85_34 ( BL34, BLN34, WL85);
sram_cell_6t_3 inst_cell_85_33 ( BL33, BLN33, WL85);
sram_cell_6t_3 inst_cell_85_32 ( BL32, BLN32, WL85);
sram_cell_6t_3 inst_cell_85_31 ( BL31, BLN31, WL85);
sram_cell_6t_3 inst_cell_85_30 ( BL30, BLN30, WL85);
sram_cell_6t_3 inst_cell_85_29 ( BL29, BLN29, WL85);
sram_cell_6t_3 inst_cell_85_28 ( BL28, BLN28, WL85);
sram_cell_6t_3 inst_cell_85_27 ( BL27, BLN27, WL85);
sram_cell_6t_3 inst_cell_85_26 ( BL26, BLN26, WL85);
sram_cell_6t_3 inst_cell_85_25 ( BL25, BLN25, WL85);
sram_cell_6t_3 inst_cell_85_24 ( BL24, BLN24, WL85);
sram_cell_6t_3 inst_cell_85_23 ( BL23, BLN23, WL85);
sram_cell_6t_3 inst_cell_85_22 ( BL22, BLN22, WL85);
sram_cell_6t_3 inst_cell_85_21 ( BL21, BLN21, WL85);
sram_cell_6t_3 inst_cell_85_20 ( BL20, BLN20, WL85);
sram_cell_6t_3 inst_cell_85_19 ( BL19, BLN19, WL85);
sram_cell_6t_3 inst_cell_85_18 ( BL18, BLN18, WL85);
sram_cell_6t_3 inst_cell_85_17 ( BL17, BLN17, WL85);
sram_cell_6t_3 inst_cell_85_16 ( BL16, BLN16, WL85);
sram_cell_6t_3 inst_cell_85_15 ( BL15, BLN15, WL85);
sram_cell_6t_3 inst_cell_85_14 ( BL14, BLN14, WL85);
sram_cell_6t_3 inst_cell_85_13 ( BL13, BLN13, WL85);
sram_cell_6t_3 inst_cell_85_12 ( BL12, BLN12, WL85);
sram_cell_6t_3 inst_cell_85_11 ( BL11, BLN11, WL85);
sram_cell_6t_3 inst_cell_85_10 ( BL10, BLN10, WL85);
sram_cell_6t_3 inst_cell_85_9 ( BL9, BLN9, WL85);
sram_cell_6t_3 inst_cell_85_8 ( BL8, BLN8, WL85);
sram_cell_6t_3 inst_cell_85_7 ( BL7, BLN7, WL85);
sram_cell_6t_3 inst_cell_85_6 ( BL6, BLN6, WL85);
sram_cell_6t_3 inst_cell_85_5 ( BL5, BLN5, WL85);
sram_cell_6t_3 inst_cell_85_4 ( BL4, BLN4, WL85);
sram_cell_6t_3 inst_cell_85_3 ( BL3, BLN3, WL85);
sram_cell_6t_3 inst_cell_85_2 ( BL2, BLN2, WL85);
sram_cell_6t_3 inst_cell_85_1 ( BL1, BLN1, WL85);
sram_cell_6t_3 inst_cell_85_0 ( BL0, BLN0, WL85);
sram_cell_6t_3 inst_cell_84_127 ( BL127, BLN127, WL84);
sram_cell_6t_3 inst_cell_84_126 ( BL126, BLN126, WL84);
sram_cell_6t_3 inst_cell_84_125 ( BL125, BLN125, WL84);
sram_cell_6t_3 inst_cell_84_124 ( BL124, BLN124, WL84);
sram_cell_6t_3 inst_cell_84_123 ( BL123, BLN123, WL84);
sram_cell_6t_3 inst_cell_84_122 ( BL122, BLN122, WL84);
sram_cell_6t_3 inst_cell_84_121 ( BL121, BLN121, WL84);
sram_cell_6t_3 inst_cell_84_120 ( BL120, BLN120, WL84);
sram_cell_6t_3 inst_cell_84_119 ( BL119, BLN119, WL84);
sram_cell_6t_3 inst_cell_84_118 ( BL118, BLN118, WL84);
sram_cell_6t_3 inst_cell_84_117 ( BL117, BLN117, WL84);
sram_cell_6t_3 inst_cell_84_116 ( BL116, BLN116, WL84);
sram_cell_6t_3 inst_cell_84_115 ( BL115, BLN115, WL84);
sram_cell_6t_3 inst_cell_84_114 ( BL114, BLN114, WL84);
sram_cell_6t_3 inst_cell_84_113 ( BL113, BLN113, WL84);
sram_cell_6t_3 inst_cell_84_112 ( BL112, BLN112, WL84);
sram_cell_6t_3 inst_cell_84_111 ( BL111, BLN111, WL84);
sram_cell_6t_3 inst_cell_84_110 ( BL110, BLN110, WL84);
sram_cell_6t_3 inst_cell_84_109 ( BL109, BLN109, WL84);
sram_cell_6t_3 inst_cell_84_108 ( BL108, BLN108, WL84);
sram_cell_6t_3 inst_cell_84_107 ( BL107, BLN107, WL84);
sram_cell_6t_3 inst_cell_84_106 ( BL106, BLN106, WL84);
sram_cell_6t_3 inst_cell_84_105 ( BL105, BLN105, WL84);
sram_cell_6t_3 inst_cell_84_104 ( BL104, BLN104, WL84);
sram_cell_6t_3 inst_cell_84_103 ( BL103, BLN103, WL84);
sram_cell_6t_3 inst_cell_84_102 ( BL102, BLN102, WL84);
sram_cell_6t_3 inst_cell_84_101 ( BL101, BLN101, WL84);
sram_cell_6t_3 inst_cell_84_100 ( BL100, BLN100, WL84);
sram_cell_6t_3 inst_cell_84_99 ( BL99, BLN99, WL84);
sram_cell_6t_3 inst_cell_84_98 ( BL98, BLN98, WL84);
sram_cell_6t_3 inst_cell_84_97 ( BL97, BLN97, WL84);
sram_cell_6t_3 inst_cell_84_96 ( BL96, BLN96, WL84);
sram_cell_6t_3 inst_cell_84_95 ( BL95, BLN95, WL84);
sram_cell_6t_3 inst_cell_84_94 ( BL94, BLN94, WL84);
sram_cell_6t_3 inst_cell_84_93 ( BL93, BLN93, WL84);
sram_cell_6t_3 inst_cell_84_92 ( BL92, BLN92, WL84);
sram_cell_6t_3 inst_cell_84_91 ( BL91, BLN91, WL84);
sram_cell_6t_3 inst_cell_84_90 ( BL90, BLN90, WL84);
sram_cell_6t_3 inst_cell_84_89 ( BL89, BLN89, WL84);
sram_cell_6t_3 inst_cell_84_88 ( BL88, BLN88, WL84);
sram_cell_6t_3 inst_cell_84_87 ( BL87, BLN87, WL84);
sram_cell_6t_3 inst_cell_84_86 ( BL86, BLN86, WL84);
sram_cell_6t_3 inst_cell_84_85 ( BL85, BLN85, WL84);
sram_cell_6t_3 inst_cell_84_84 ( BL84, BLN84, WL84);
sram_cell_6t_3 inst_cell_84_83 ( BL83, BLN83, WL84);
sram_cell_6t_3 inst_cell_84_82 ( BL82, BLN82, WL84);
sram_cell_6t_3 inst_cell_84_81 ( BL81, BLN81, WL84);
sram_cell_6t_3 inst_cell_84_80 ( BL80, BLN80, WL84);
sram_cell_6t_3 inst_cell_84_79 ( BL79, BLN79, WL84);
sram_cell_6t_3 inst_cell_84_78 ( BL78, BLN78, WL84);
sram_cell_6t_3 inst_cell_84_77 ( BL77, BLN77, WL84);
sram_cell_6t_3 inst_cell_84_76 ( BL76, BLN76, WL84);
sram_cell_6t_3 inst_cell_84_75 ( BL75, BLN75, WL84);
sram_cell_6t_3 inst_cell_84_74 ( BL74, BLN74, WL84);
sram_cell_6t_3 inst_cell_84_73 ( BL73, BLN73, WL84);
sram_cell_6t_3 inst_cell_84_72 ( BL72, BLN72, WL84);
sram_cell_6t_3 inst_cell_84_71 ( BL71, BLN71, WL84);
sram_cell_6t_3 inst_cell_84_70 ( BL70, BLN70, WL84);
sram_cell_6t_3 inst_cell_84_69 ( BL69, BLN69, WL84);
sram_cell_6t_3 inst_cell_84_68 ( BL68, BLN68, WL84);
sram_cell_6t_3 inst_cell_84_67 ( BL67, BLN67, WL84);
sram_cell_6t_3 inst_cell_84_66 ( BL66, BLN66, WL84);
sram_cell_6t_3 inst_cell_84_65 ( BL65, BLN65, WL84);
sram_cell_6t_3 inst_cell_84_64 ( BL64, BLN64, WL84);
sram_cell_6t_3 inst_cell_84_63 ( BL63, BLN63, WL84);
sram_cell_6t_3 inst_cell_84_62 ( BL62, BLN62, WL84);
sram_cell_6t_3 inst_cell_84_61 ( BL61, BLN61, WL84);
sram_cell_6t_3 inst_cell_84_60 ( BL60, BLN60, WL84);
sram_cell_6t_3 inst_cell_84_59 ( BL59, BLN59, WL84);
sram_cell_6t_3 inst_cell_84_58 ( BL58, BLN58, WL84);
sram_cell_6t_3 inst_cell_84_57 ( BL57, BLN57, WL84);
sram_cell_6t_3 inst_cell_84_56 ( BL56, BLN56, WL84);
sram_cell_6t_3 inst_cell_84_55 ( BL55, BLN55, WL84);
sram_cell_6t_3 inst_cell_84_54 ( BL54, BLN54, WL84);
sram_cell_6t_3 inst_cell_84_53 ( BL53, BLN53, WL84);
sram_cell_6t_3 inst_cell_84_52 ( BL52, BLN52, WL84);
sram_cell_6t_3 inst_cell_84_51 ( BL51, BLN51, WL84);
sram_cell_6t_3 inst_cell_84_50 ( BL50, BLN50, WL84);
sram_cell_6t_3 inst_cell_84_49 ( BL49, BLN49, WL84);
sram_cell_6t_3 inst_cell_84_48 ( BL48, BLN48, WL84);
sram_cell_6t_3 inst_cell_84_47 ( BL47, BLN47, WL84);
sram_cell_6t_3 inst_cell_84_46 ( BL46, BLN46, WL84);
sram_cell_6t_3 inst_cell_84_45 ( BL45, BLN45, WL84);
sram_cell_6t_3 inst_cell_84_44 ( BL44, BLN44, WL84);
sram_cell_6t_3 inst_cell_84_43 ( BL43, BLN43, WL84);
sram_cell_6t_3 inst_cell_84_42 ( BL42, BLN42, WL84);
sram_cell_6t_3 inst_cell_84_41 ( BL41, BLN41, WL84);
sram_cell_6t_3 inst_cell_84_40 ( BL40, BLN40, WL84);
sram_cell_6t_3 inst_cell_84_39 ( BL39, BLN39, WL84);
sram_cell_6t_3 inst_cell_84_38 ( BL38, BLN38, WL84);
sram_cell_6t_3 inst_cell_84_37 ( BL37, BLN37, WL84);
sram_cell_6t_3 inst_cell_84_36 ( BL36, BLN36, WL84);
sram_cell_6t_3 inst_cell_84_35 ( BL35, BLN35, WL84);
sram_cell_6t_3 inst_cell_84_34 ( BL34, BLN34, WL84);
sram_cell_6t_3 inst_cell_84_33 ( BL33, BLN33, WL84);
sram_cell_6t_3 inst_cell_84_32 ( BL32, BLN32, WL84);
sram_cell_6t_3 inst_cell_84_31 ( BL31, BLN31, WL84);
sram_cell_6t_3 inst_cell_84_30 ( BL30, BLN30, WL84);
sram_cell_6t_3 inst_cell_84_29 ( BL29, BLN29, WL84);
sram_cell_6t_3 inst_cell_84_28 ( BL28, BLN28, WL84);
sram_cell_6t_3 inst_cell_84_27 ( BL27, BLN27, WL84);
sram_cell_6t_3 inst_cell_84_26 ( BL26, BLN26, WL84);
sram_cell_6t_3 inst_cell_84_25 ( BL25, BLN25, WL84);
sram_cell_6t_3 inst_cell_84_24 ( BL24, BLN24, WL84);
sram_cell_6t_3 inst_cell_84_23 ( BL23, BLN23, WL84);
sram_cell_6t_3 inst_cell_84_22 ( BL22, BLN22, WL84);
sram_cell_6t_3 inst_cell_84_21 ( BL21, BLN21, WL84);
sram_cell_6t_3 inst_cell_84_20 ( BL20, BLN20, WL84);
sram_cell_6t_3 inst_cell_84_19 ( BL19, BLN19, WL84);
sram_cell_6t_3 inst_cell_84_18 ( BL18, BLN18, WL84);
sram_cell_6t_3 inst_cell_84_17 ( BL17, BLN17, WL84);
sram_cell_6t_3 inst_cell_84_16 ( BL16, BLN16, WL84);
sram_cell_6t_3 inst_cell_84_15 ( BL15, BLN15, WL84);
sram_cell_6t_3 inst_cell_84_14 ( BL14, BLN14, WL84);
sram_cell_6t_3 inst_cell_84_13 ( BL13, BLN13, WL84);
sram_cell_6t_3 inst_cell_84_12 ( BL12, BLN12, WL84);
sram_cell_6t_3 inst_cell_84_11 ( BL11, BLN11, WL84);
sram_cell_6t_3 inst_cell_84_10 ( BL10, BLN10, WL84);
sram_cell_6t_3 inst_cell_84_9 ( BL9, BLN9, WL84);
sram_cell_6t_3 inst_cell_84_8 ( BL8, BLN8, WL84);
sram_cell_6t_3 inst_cell_84_7 ( BL7, BLN7, WL84);
sram_cell_6t_3 inst_cell_84_6 ( BL6, BLN6, WL84);
sram_cell_6t_3 inst_cell_84_5 ( BL5, BLN5, WL84);
sram_cell_6t_3 inst_cell_84_4 ( BL4, BLN4, WL84);
sram_cell_6t_3 inst_cell_84_3 ( BL3, BLN3, WL84);
sram_cell_6t_3 inst_cell_84_2 ( BL2, BLN2, WL84);
sram_cell_6t_3 inst_cell_84_1 ( BL1, BLN1, WL84);
sram_cell_6t_3 inst_cell_84_0 ( BL0, BLN0, WL84);
sram_cell_6t_3 inst_cell_83_127 ( BL127, BLN127, WL83);
sram_cell_6t_3 inst_cell_83_126 ( BL126, BLN126, WL83);
sram_cell_6t_3 inst_cell_83_125 ( BL125, BLN125, WL83);
sram_cell_6t_3 inst_cell_83_124 ( BL124, BLN124, WL83);
sram_cell_6t_3 inst_cell_83_123 ( BL123, BLN123, WL83);
sram_cell_6t_3 inst_cell_83_122 ( BL122, BLN122, WL83);
sram_cell_6t_3 inst_cell_83_121 ( BL121, BLN121, WL83);
sram_cell_6t_3 inst_cell_83_120 ( BL120, BLN120, WL83);
sram_cell_6t_3 inst_cell_83_119 ( BL119, BLN119, WL83);
sram_cell_6t_3 inst_cell_83_118 ( BL118, BLN118, WL83);
sram_cell_6t_3 inst_cell_83_117 ( BL117, BLN117, WL83);
sram_cell_6t_3 inst_cell_83_116 ( BL116, BLN116, WL83);
sram_cell_6t_3 inst_cell_83_115 ( BL115, BLN115, WL83);
sram_cell_6t_3 inst_cell_83_114 ( BL114, BLN114, WL83);
sram_cell_6t_3 inst_cell_83_113 ( BL113, BLN113, WL83);
sram_cell_6t_3 inst_cell_83_112 ( BL112, BLN112, WL83);
sram_cell_6t_3 inst_cell_83_111 ( BL111, BLN111, WL83);
sram_cell_6t_3 inst_cell_83_110 ( BL110, BLN110, WL83);
sram_cell_6t_3 inst_cell_83_109 ( BL109, BLN109, WL83);
sram_cell_6t_3 inst_cell_83_108 ( BL108, BLN108, WL83);
sram_cell_6t_3 inst_cell_83_107 ( BL107, BLN107, WL83);
sram_cell_6t_3 inst_cell_83_106 ( BL106, BLN106, WL83);
sram_cell_6t_3 inst_cell_83_105 ( BL105, BLN105, WL83);
sram_cell_6t_3 inst_cell_83_104 ( BL104, BLN104, WL83);
sram_cell_6t_3 inst_cell_83_103 ( BL103, BLN103, WL83);
sram_cell_6t_3 inst_cell_83_102 ( BL102, BLN102, WL83);
sram_cell_6t_3 inst_cell_83_101 ( BL101, BLN101, WL83);
sram_cell_6t_3 inst_cell_83_100 ( BL100, BLN100, WL83);
sram_cell_6t_3 inst_cell_83_99 ( BL99, BLN99, WL83);
sram_cell_6t_3 inst_cell_83_98 ( BL98, BLN98, WL83);
sram_cell_6t_3 inst_cell_83_97 ( BL97, BLN97, WL83);
sram_cell_6t_3 inst_cell_83_96 ( BL96, BLN96, WL83);
sram_cell_6t_3 inst_cell_83_95 ( BL95, BLN95, WL83);
sram_cell_6t_3 inst_cell_83_94 ( BL94, BLN94, WL83);
sram_cell_6t_3 inst_cell_83_93 ( BL93, BLN93, WL83);
sram_cell_6t_3 inst_cell_83_92 ( BL92, BLN92, WL83);
sram_cell_6t_3 inst_cell_83_91 ( BL91, BLN91, WL83);
sram_cell_6t_3 inst_cell_83_90 ( BL90, BLN90, WL83);
sram_cell_6t_3 inst_cell_83_89 ( BL89, BLN89, WL83);
sram_cell_6t_3 inst_cell_83_88 ( BL88, BLN88, WL83);
sram_cell_6t_3 inst_cell_83_87 ( BL87, BLN87, WL83);
sram_cell_6t_3 inst_cell_83_86 ( BL86, BLN86, WL83);
sram_cell_6t_3 inst_cell_83_85 ( BL85, BLN85, WL83);
sram_cell_6t_3 inst_cell_83_84 ( BL84, BLN84, WL83);
sram_cell_6t_3 inst_cell_83_83 ( BL83, BLN83, WL83);
sram_cell_6t_3 inst_cell_83_82 ( BL82, BLN82, WL83);
sram_cell_6t_3 inst_cell_83_81 ( BL81, BLN81, WL83);
sram_cell_6t_3 inst_cell_83_80 ( BL80, BLN80, WL83);
sram_cell_6t_3 inst_cell_83_79 ( BL79, BLN79, WL83);
sram_cell_6t_3 inst_cell_83_78 ( BL78, BLN78, WL83);
sram_cell_6t_3 inst_cell_83_77 ( BL77, BLN77, WL83);
sram_cell_6t_3 inst_cell_83_76 ( BL76, BLN76, WL83);
sram_cell_6t_3 inst_cell_83_75 ( BL75, BLN75, WL83);
sram_cell_6t_3 inst_cell_83_74 ( BL74, BLN74, WL83);
sram_cell_6t_3 inst_cell_83_73 ( BL73, BLN73, WL83);
sram_cell_6t_3 inst_cell_83_72 ( BL72, BLN72, WL83);
sram_cell_6t_3 inst_cell_83_71 ( BL71, BLN71, WL83);
sram_cell_6t_3 inst_cell_83_70 ( BL70, BLN70, WL83);
sram_cell_6t_3 inst_cell_83_69 ( BL69, BLN69, WL83);
sram_cell_6t_3 inst_cell_83_68 ( BL68, BLN68, WL83);
sram_cell_6t_3 inst_cell_83_67 ( BL67, BLN67, WL83);
sram_cell_6t_3 inst_cell_83_66 ( BL66, BLN66, WL83);
sram_cell_6t_3 inst_cell_83_65 ( BL65, BLN65, WL83);
sram_cell_6t_3 inst_cell_83_64 ( BL64, BLN64, WL83);
sram_cell_6t_3 inst_cell_83_63 ( BL63, BLN63, WL83);
sram_cell_6t_3 inst_cell_83_62 ( BL62, BLN62, WL83);
sram_cell_6t_3 inst_cell_83_61 ( BL61, BLN61, WL83);
sram_cell_6t_3 inst_cell_83_60 ( BL60, BLN60, WL83);
sram_cell_6t_3 inst_cell_83_59 ( BL59, BLN59, WL83);
sram_cell_6t_3 inst_cell_83_58 ( BL58, BLN58, WL83);
sram_cell_6t_3 inst_cell_83_57 ( BL57, BLN57, WL83);
sram_cell_6t_3 inst_cell_83_56 ( BL56, BLN56, WL83);
sram_cell_6t_3 inst_cell_83_55 ( BL55, BLN55, WL83);
sram_cell_6t_3 inst_cell_83_54 ( BL54, BLN54, WL83);
sram_cell_6t_3 inst_cell_83_53 ( BL53, BLN53, WL83);
sram_cell_6t_3 inst_cell_83_52 ( BL52, BLN52, WL83);
sram_cell_6t_3 inst_cell_83_51 ( BL51, BLN51, WL83);
sram_cell_6t_3 inst_cell_83_50 ( BL50, BLN50, WL83);
sram_cell_6t_3 inst_cell_83_49 ( BL49, BLN49, WL83);
sram_cell_6t_3 inst_cell_83_48 ( BL48, BLN48, WL83);
sram_cell_6t_3 inst_cell_83_47 ( BL47, BLN47, WL83);
sram_cell_6t_3 inst_cell_83_46 ( BL46, BLN46, WL83);
sram_cell_6t_3 inst_cell_83_45 ( BL45, BLN45, WL83);
sram_cell_6t_3 inst_cell_83_44 ( BL44, BLN44, WL83);
sram_cell_6t_3 inst_cell_83_43 ( BL43, BLN43, WL83);
sram_cell_6t_3 inst_cell_83_42 ( BL42, BLN42, WL83);
sram_cell_6t_3 inst_cell_83_41 ( BL41, BLN41, WL83);
sram_cell_6t_3 inst_cell_83_40 ( BL40, BLN40, WL83);
sram_cell_6t_3 inst_cell_83_39 ( BL39, BLN39, WL83);
sram_cell_6t_3 inst_cell_83_38 ( BL38, BLN38, WL83);
sram_cell_6t_3 inst_cell_83_37 ( BL37, BLN37, WL83);
sram_cell_6t_3 inst_cell_83_36 ( BL36, BLN36, WL83);
sram_cell_6t_3 inst_cell_83_35 ( BL35, BLN35, WL83);
sram_cell_6t_3 inst_cell_83_34 ( BL34, BLN34, WL83);
sram_cell_6t_3 inst_cell_83_33 ( BL33, BLN33, WL83);
sram_cell_6t_3 inst_cell_83_32 ( BL32, BLN32, WL83);
sram_cell_6t_3 inst_cell_83_31 ( BL31, BLN31, WL83);
sram_cell_6t_3 inst_cell_83_30 ( BL30, BLN30, WL83);
sram_cell_6t_3 inst_cell_83_29 ( BL29, BLN29, WL83);
sram_cell_6t_3 inst_cell_83_28 ( BL28, BLN28, WL83);
sram_cell_6t_3 inst_cell_83_27 ( BL27, BLN27, WL83);
sram_cell_6t_3 inst_cell_83_26 ( BL26, BLN26, WL83);
sram_cell_6t_3 inst_cell_83_25 ( BL25, BLN25, WL83);
sram_cell_6t_3 inst_cell_83_24 ( BL24, BLN24, WL83);
sram_cell_6t_3 inst_cell_83_23 ( BL23, BLN23, WL83);
sram_cell_6t_3 inst_cell_83_22 ( BL22, BLN22, WL83);
sram_cell_6t_3 inst_cell_83_21 ( BL21, BLN21, WL83);
sram_cell_6t_3 inst_cell_83_20 ( BL20, BLN20, WL83);
sram_cell_6t_3 inst_cell_83_19 ( BL19, BLN19, WL83);
sram_cell_6t_3 inst_cell_83_18 ( BL18, BLN18, WL83);
sram_cell_6t_3 inst_cell_83_17 ( BL17, BLN17, WL83);
sram_cell_6t_3 inst_cell_83_16 ( BL16, BLN16, WL83);
sram_cell_6t_3 inst_cell_83_15 ( BL15, BLN15, WL83);
sram_cell_6t_3 inst_cell_83_14 ( BL14, BLN14, WL83);
sram_cell_6t_3 inst_cell_83_13 ( BL13, BLN13, WL83);
sram_cell_6t_3 inst_cell_83_12 ( BL12, BLN12, WL83);
sram_cell_6t_3 inst_cell_83_11 ( BL11, BLN11, WL83);
sram_cell_6t_3 inst_cell_83_10 ( BL10, BLN10, WL83);
sram_cell_6t_3 inst_cell_83_9 ( BL9, BLN9, WL83);
sram_cell_6t_3 inst_cell_83_8 ( BL8, BLN8, WL83);
sram_cell_6t_3 inst_cell_83_7 ( BL7, BLN7, WL83);
sram_cell_6t_3 inst_cell_83_6 ( BL6, BLN6, WL83);
sram_cell_6t_3 inst_cell_83_5 ( BL5, BLN5, WL83);
sram_cell_6t_3 inst_cell_83_4 ( BL4, BLN4, WL83);
sram_cell_6t_3 inst_cell_83_3 ( BL3, BLN3, WL83);
sram_cell_6t_3 inst_cell_83_2 ( BL2, BLN2, WL83);
sram_cell_6t_3 inst_cell_83_1 ( BL1, BLN1, WL83);
sram_cell_6t_3 inst_cell_83_0 ( BL0, BLN0, WL83);
sram_cell_6t_3 inst_cell_82_127 ( BL127, BLN127, WL82);
sram_cell_6t_3 inst_cell_82_126 ( BL126, BLN126, WL82);
sram_cell_6t_3 inst_cell_82_125 ( BL125, BLN125, WL82);
sram_cell_6t_3 inst_cell_82_124 ( BL124, BLN124, WL82);
sram_cell_6t_3 inst_cell_82_123 ( BL123, BLN123, WL82);
sram_cell_6t_3 inst_cell_82_122 ( BL122, BLN122, WL82);
sram_cell_6t_3 inst_cell_82_121 ( BL121, BLN121, WL82);
sram_cell_6t_3 inst_cell_82_120 ( BL120, BLN120, WL82);
sram_cell_6t_3 inst_cell_82_119 ( BL119, BLN119, WL82);
sram_cell_6t_3 inst_cell_82_118 ( BL118, BLN118, WL82);
sram_cell_6t_3 inst_cell_82_117 ( BL117, BLN117, WL82);
sram_cell_6t_3 inst_cell_82_116 ( BL116, BLN116, WL82);
sram_cell_6t_3 inst_cell_82_115 ( BL115, BLN115, WL82);
sram_cell_6t_3 inst_cell_82_114 ( BL114, BLN114, WL82);
sram_cell_6t_3 inst_cell_82_113 ( BL113, BLN113, WL82);
sram_cell_6t_3 inst_cell_82_112 ( BL112, BLN112, WL82);
sram_cell_6t_3 inst_cell_82_111 ( BL111, BLN111, WL82);
sram_cell_6t_3 inst_cell_82_110 ( BL110, BLN110, WL82);
sram_cell_6t_3 inst_cell_82_109 ( BL109, BLN109, WL82);
sram_cell_6t_3 inst_cell_82_108 ( BL108, BLN108, WL82);
sram_cell_6t_3 inst_cell_82_107 ( BL107, BLN107, WL82);
sram_cell_6t_3 inst_cell_82_106 ( BL106, BLN106, WL82);
sram_cell_6t_3 inst_cell_82_105 ( BL105, BLN105, WL82);
sram_cell_6t_3 inst_cell_82_104 ( BL104, BLN104, WL82);
sram_cell_6t_3 inst_cell_82_103 ( BL103, BLN103, WL82);
sram_cell_6t_3 inst_cell_82_102 ( BL102, BLN102, WL82);
sram_cell_6t_3 inst_cell_82_101 ( BL101, BLN101, WL82);
sram_cell_6t_3 inst_cell_82_100 ( BL100, BLN100, WL82);
sram_cell_6t_3 inst_cell_82_99 ( BL99, BLN99, WL82);
sram_cell_6t_3 inst_cell_82_98 ( BL98, BLN98, WL82);
sram_cell_6t_3 inst_cell_82_97 ( BL97, BLN97, WL82);
sram_cell_6t_3 inst_cell_82_96 ( BL96, BLN96, WL82);
sram_cell_6t_3 inst_cell_82_95 ( BL95, BLN95, WL82);
sram_cell_6t_3 inst_cell_82_94 ( BL94, BLN94, WL82);
sram_cell_6t_3 inst_cell_82_93 ( BL93, BLN93, WL82);
sram_cell_6t_3 inst_cell_82_92 ( BL92, BLN92, WL82);
sram_cell_6t_3 inst_cell_82_91 ( BL91, BLN91, WL82);
sram_cell_6t_3 inst_cell_82_90 ( BL90, BLN90, WL82);
sram_cell_6t_3 inst_cell_82_89 ( BL89, BLN89, WL82);
sram_cell_6t_3 inst_cell_82_88 ( BL88, BLN88, WL82);
sram_cell_6t_3 inst_cell_82_87 ( BL87, BLN87, WL82);
sram_cell_6t_3 inst_cell_82_86 ( BL86, BLN86, WL82);
sram_cell_6t_3 inst_cell_82_85 ( BL85, BLN85, WL82);
sram_cell_6t_3 inst_cell_82_84 ( BL84, BLN84, WL82);
sram_cell_6t_3 inst_cell_82_83 ( BL83, BLN83, WL82);
sram_cell_6t_3 inst_cell_82_82 ( BL82, BLN82, WL82);
sram_cell_6t_3 inst_cell_82_81 ( BL81, BLN81, WL82);
sram_cell_6t_3 inst_cell_82_80 ( BL80, BLN80, WL82);
sram_cell_6t_3 inst_cell_82_79 ( BL79, BLN79, WL82);
sram_cell_6t_3 inst_cell_82_78 ( BL78, BLN78, WL82);
sram_cell_6t_3 inst_cell_82_77 ( BL77, BLN77, WL82);
sram_cell_6t_3 inst_cell_82_76 ( BL76, BLN76, WL82);
sram_cell_6t_3 inst_cell_82_75 ( BL75, BLN75, WL82);
sram_cell_6t_3 inst_cell_82_74 ( BL74, BLN74, WL82);
sram_cell_6t_3 inst_cell_82_73 ( BL73, BLN73, WL82);
sram_cell_6t_3 inst_cell_82_72 ( BL72, BLN72, WL82);
sram_cell_6t_3 inst_cell_82_71 ( BL71, BLN71, WL82);
sram_cell_6t_3 inst_cell_82_70 ( BL70, BLN70, WL82);
sram_cell_6t_3 inst_cell_82_69 ( BL69, BLN69, WL82);
sram_cell_6t_3 inst_cell_82_68 ( BL68, BLN68, WL82);
sram_cell_6t_3 inst_cell_82_67 ( BL67, BLN67, WL82);
sram_cell_6t_3 inst_cell_82_66 ( BL66, BLN66, WL82);
sram_cell_6t_3 inst_cell_82_65 ( BL65, BLN65, WL82);
sram_cell_6t_3 inst_cell_82_64 ( BL64, BLN64, WL82);
sram_cell_6t_3 inst_cell_82_63 ( BL63, BLN63, WL82);
sram_cell_6t_3 inst_cell_82_62 ( BL62, BLN62, WL82);
sram_cell_6t_3 inst_cell_82_61 ( BL61, BLN61, WL82);
sram_cell_6t_3 inst_cell_82_60 ( BL60, BLN60, WL82);
sram_cell_6t_3 inst_cell_82_59 ( BL59, BLN59, WL82);
sram_cell_6t_3 inst_cell_82_58 ( BL58, BLN58, WL82);
sram_cell_6t_3 inst_cell_82_57 ( BL57, BLN57, WL82);
sram_cell_6t_3 inst_cell_82_56 ( BL56, BLN56, WL82);
sram_cell_6t_3 inst_cell_82_55 ( BL55, BLN55, WL82);
sram_cell_6t_3 inst_cell_82_54 ( BL54, BLN54, WL82);
sram_cell_6t_3 inst_cell_82_53 ( BL53, BLN53, WL82);
sram_cell_6t_3 inst_cell_82_52 ( BL52, BLN52, WL82);
sram_cell_6t_3 inst_cell_82_51 ( BL51, BLN51, WL82);
sram_cell_6t_3 inst_cell_82_50 ( BL50, BLN50, WL82);
sram_cell_6t_3 inst_cell_82_49 ( BL49, BLN49, WL82);
sram_cell_6t_3 inst_cell_82_48 ( BL48, BLN48, WL82);
sram_cell_6t_3 inst_cell_82_47 ( BL47, BLN47, WL82);
sram_cell_6t_3 inst_cell_82_46 ( BL46, BLN46, WL82);
sram_cell_6t_3 inst_cell_82_45 ( BL45, BLN45, WL82);
sram_cell_6t_3 inst_cell_82_44 ( BL44, BLN44, WL82);
sram_cell_6t_3 inst_cell_82_43 ( BL43, BLN43, WL82);
sram_cell_6t_3 inst_cell_82_42 ( BL42, BLN42, WL82);
sram_cell_6t_3 inst_cell_82_41 ( BL41, BLN41, WL82);
sram_cell_6t_3 inst_cell_82_40 ( BL40, BLN40, WL82);
sram_cell_6t_3 inst_cell_82_39 ( BL39, BLN39, WL82);
sram_cell_6t_3 inst_cell_82_38 ( BL38, BLN38, WL82);
sram_cell_6t_3 inst_cell_82_37 ( BL37, BLN37, WL82);
sram_cell_6t_3 inst_cell_82_36 ( BL36, BLN36, WL82);
sram_cell_6t_3 inst_cell_82_35 ( BL35, BLN35, WL82);
sram_cell_6t_3 inst_cell_82_34 ( BL34, BLN34, WL82);
sram_cell_6t_3 inst_cell_82_33 ( BL33, BLN33, WL82);
sram_cell_6t_3 inst_cell_82_32 ( BL32, BLN32, WL82);
sram_cell_6t_3 inst_cell_82_31 ( BL31, BLN31, WL82);
sram_cell_6t_3 inst_cell_82_30 ( BL30, BLN30, WL82);
sram_cell_6t_3 inst_cell_82_29 ( BL29, BLN29, WL82);
sram_cell_6t_3 inst_cell_82_28 ( BL28, BLN28, WL82);
sram_cell_6t_3 inst_cell_82_27 ( BL27, BLN27, WL82);
sram_cell_6t_3 inst_cell_82_26 ( BL26, BLN26, WL82);
sram_cell_6t_3 inst_cell_82_25 ( BL25, BLN25, WL82);
sram_cell_6t_3 inst_cell_82_24 ( BL24, BLN24, WL82);
sram_cell_6t_3 inst_cell_82_23 ( BL23, BLN23, WL82);
sram_cell_6t_3 inst_cell_82_22 ( BL22, BLN22, WL82);
sram_cell_6t_3 inst_cell_82_21 ( BL21, BLN21, WL82);
sram_cell_6t_3 inst_cell_82_20 ( BL20, BLN20, WL82);
sram_cell_6t_3 inst_cell_82_19 ( BL19, BLN19, WL82);
sram_cell_6t_3 inst_cell_82_18 ( BL18, BLN18, WL82);
sram_cell_6t_3 inst_cell_82_17 ( BL17, BLN17, WL82);
sram_cell_6t_3 inst_cell_82_16 ( BL16, BLN16, WL82);
sram_cell_6t_3 inst_cell_82_15 ( BL15, BLN15, WL82);
sram_cell_6t_3 inst_cell_82_14 ( BL14, BLN14, WL82);
sram_cell_6t_3 inst_cell_82_13 ( BL13, BLN13, WL82);
sram_cell_6t_3 inst_cell_82_12 ( BL12, BLN12, WL82);
sram_cell_6t_3 inst_cell_82_11 ( BL11, BLN11, WL82);
sram_cell_6t_3 inst_cell_82_10 ( BL10, BLN10, WL82);
sram_cell_6t_3 inst_cell_82_9 ( BL9, BLN9, WL82);
sram_cell_6t_3 inst_cell_82_8 ( BL8, BLN8, WL82);
sram_cell_6t_3 inst_cell_82_7 ( BL7, BLN7, WL82);
sram_cell_6t_3 inst_cell_82_6 ( BL6, BLN6, WL82);
sram_cell_6t_3 inst_cell_82_5 ( BL5, BLN5, WL82);
sram_cell_6t_3 inst_cell_82_4 ( BL4, BLN4, WL82);
sram_cell_6t_3 inst_cell_82_3 ( BL3, BLN3, WL82);
sram_cell_6t_3 inst_cell_82_2 ( BL2, BLN2, WL82);
sram_cell_6t_3 inst_cell_82_1 ( BL1, BLN1, WL82);
sram_cell_6t_3 inst_cell_82_0 ( BL0, BLN0, WL82);
sram_cell_6t_3 inst_cell_81_127 ( BL127, BLN127, WL81);
sram_cell_6t_3 inst_cell_81_126 ( BL126, BLN126, WL81);
sram_cell_6t_3 inst_cell_81_125 ( BL125, BLN125, WL81);
sram_cell_6t_3 inst_cell_81_124 ( BL124, BLN124, WL81);
sram_cell_6t_3 inst_cell_81_123 ( BL123, BLN123, WL81);
sram_cell_6t_3 inst_cell_81_122 ( BL122, BLN122, WL81);
sram_cell_6t_3 inst_cell_81_121 ( BL121, BLN121, WL81);
sram_cell_6t_3 inst_cell_81_120 ( BL120, BLN120, WL81);
sram_cell_6t_3 inst_cell_81_119 ( BL119, BLN119, WL81);
sram_cell_6t_3 inst_cell_81_118 ( BL118, BLN118, WL81);
sram_cell_6t_3 inst_cell_81_117 ( BL117, BLN117, WL81);
sram_cell_6t_3 inst_cell_81_116 ( BL116, BLN116, WL81);
sram_cell_6t_3 inst_cell_81_115 ( BL115, BLN115, WL81);
sram_cell_6t_3 inst_cell_81_114 ( BL114, BLN114, WL81);
sram_cell_6t_3 inst_cell_81_113 ( BL113, BLN113, WL81);
sram_cell_6t_3 inst_cell_81_112 ( BL112, BLN112, WL81);
sram_cell_6t_3 inst_cell_81_111 ( BL111, BLN111, WL81);
sram_cell_6t_3 inst_cell_81_110 ( BL110, BLN110, WL81);
sram_cell_6t_3 inst_cell_81_109 ( BL109, BLN109, WL81);
sram_cell_6t_3 inst_cell_81_108 ( BL108, BLN108, WL81);
sram_cell_6t_3 inst_cell_81_107 ( BL107, BLN107, WL81);
sram_cell_6t_3 inst_cell_81_106 ( BL106, BLN106, WL81);
sram_cell_6t_3 inst_cell_81_105 ( BL105, BLN105, WL81);
sram_cell_6t_3 inst_cell_81_104 ( BL104, BLN104, WL81);
sram_cell_6t_3 inst_cell_81_103 ( BL103, BLN103, WL81);
sram_cell_6t_3 inst_cell_81_102 ( BL102, BLN102, WL81);
sram_cell_6t_3 inst_cell_81_101 ( BL101, BLN101, WL81);
sram_cell_6t_3 inst_cell_81_100 ( BL100, BLN100, WL81);
sram_cell_6t_3 inst_cell_81_99 ( BL99, BLN99, WL81);
sram_cell_6t_3 inst_cell_81_98 ( BL98, BLN98, WL81);
sram_cell_6t_3 inst_cell_81_97 ( BL97, BLN97, WL81);
sram_cell_6t_3 inst_cell_81_96 ( BL96, BLN96, WL81);
sram_cell_6t_3 inst_cell_81_95 ( BL95, BLN95, WL81);
sram_cell_6t_3 inst_cell_81_94 ( BL94, BLN94, WL81);
sram_cell_6t_3 inst_cell_81_93 ( BL93, BLN93, WL81);
sram_cell_6t_3 inst_cell_81_92 ( BL92, BLN92, WL81);
sram_cell_6t_3 inst_cell_81_91 ( BL91, BLN91, WL81);
sram_cell_6t_3 inst_cell_81_90 ( BL90, BLN90, WL81);
sram_cell_6t_3 inst_cell_81_89 ( BL89, BLN89, WL81);
sram_cell_6t_3 inst_cell_81_88 ( BL88, BLN88, WL81);
sram_cell_6t_3 inst_cell_81_87 ( BL87, BLN87, WL81);
sram_cell_6t_3 inst_cell_81_86 ( BL86, BLN86, WL81);
sram_cell_6t_3 inst_cell_81_85 ( BL85, BLN85, WL81);
sram_cell_6t_3 inst_cell_81_84 ( BL84, BLN84, WL81);
sram_cell_6t_3 inst_cell_81_83 ( BL83, BLN83, WL81);
sram_cell_6t_3 inst_cell_81_82 ( BL82, BLN82, WL81);
sram_cell_6t_3 inst_cell_81_81 ( BL81, BLN81, WL81);
sram_cell_6t_3 inst_cell_81_80 ( BL80, BLN80, WL81);
sram_cell_6t_3 inst_cell_81_79 ( BL79, BLN79, WL81);
sram_cell_6t_3 inst_cell_81_78 ( BL78, BLN78, WL81);
sram_cell_6t_3 inst_cell_81_77 ( BL77, BLN77, WL81);
sram_cell_6t_3 inst_cell_81_76 ( BL76, BLN76, WL81);
sram_cell_6t_3 inst_cell_81_75 ( BL75, BLN75, WL81);
sram_cell_6t_3 inst_cell_81_74 ( BL74, BLN74, WL81);
sram_cell_6t_3 inst_cell_81_73 ( BL73, BLN73, WL81);
sram_cell_6t_3 inst_cell_81_72 ( BL72, BLN72, WL81);
sram_cell_6t_3 inst_cell_81_71 ( BL71, BLN71, WL81);
sram_cell_6t_3 inst_cell_81_70 ( BL70, BLN70, WL81);
sram_cell_6t_3 inst_cell_81_69 ( BL69, BLN69, WL81);
sram_cell_6t_3 inst_cell_81_68 ( BL68, BLN68, WL81);
sram_cell_6t_3 inst_cell_81_67 ( BL67, BLN67, WL81);
sram_cell_6t_3 inst_cell_81_66 ( BL66, BLN66, WL81);
sram_cell_6t_3 inst_cell_81_65 ( BL65, BLN65, WL81);
sram_cell_6t_3 inst_cell_81_64 ( BL64, BLN64, WL81);
sram_cell_6t_3 inst_cell_81_63 ( BL63, BLN63, WL81);
sram_cell_6t_3 inst_cell_81_62 ( BL62, BLN62, WL81);
sram_cell_6t_3 inst_cell_81_61 ( BL61, BLN61, WL81);
sram_cell_6t_3 inst_cell_81_60 ( BL60, BLN60, WL81);
sram_cell_6t_3 inst_cell_81_59 ( BL59, BLN59, WL81);
sram_cell_6t_3 inst_cell_81_58 ( BL58, BLN58, WL81);
sram_cell_6t_3 inst_cell_81_57 ( BL57, BLN57, WL81);
sram_cell_6t_3 inst_cell_81_56 ( BL56, BLN56, WL81);
sram_cell_6t_3 inst_cell_81_55 ( BL55, BLN55, WL81);
sram_cell_6t_3 inst_cell_81_54 ( BL54, BLN54, WL81);
sram_cell_6t_3 inst_cell_81_53 ( BL53, BLN53, WL81);
sram_cell_6t_3 inst_cell_81_52 ( BL52, BLN52, WL81);
sram_cell_6t_3 inst_cell_81_51 ( BL51, BLN51, WL81);
sram_cell_6t_3 inst_cell_81_50 ( BL50, BLN50, WL81);
sram_cell_6t_3 inst_cell_81_49 ( BL49, BLN49, WL81);
sram_cell_6t_3 inst_cell_81_48 ( BL48, BLN48, WL81);
sram_cell_6t_3 inst_cell_81_47 ( BL47, BLN47, WL81);
sram_cell_6t_3 inst_cell_81_46 ( BL46, BLN46, WL81);
sram_cell_6t_3 inst_cell_81_45 ( BL45, BLN45, WL81);
sram_cell_6t_3 inst_cell_81_44 ( BL44, BLN44, WL81);
sram_cell_6t_3 inst_cell_81_43 ( BL43, BLN43, WL81);
sram_cell_6t_3 inst_cell_81_42 ( BL42, BLN42, WL81);
sram_cell_6t_3 inst_cell_81_41 ( BL41, BLN41, WL81);
sram_cell_6t_3 inst_cell_81_40 ( BL40, BLN40, WL81);
sram_cell_6t_3 inst_cell_81_39 ( BL39, BLN39, WL81);
sram_cell_6t_3 inst_cell_81_38 ( BL38, BLN38, WL81);
sram_cell_6t_3 inst_cell_81_37 ( BL37, BLN37, WL81);
sram_cell_6t_3 inst_cell_81_36 ( BL36, BLN36, WL81);
sram_cell_6t_3 inst_cell_81_35 ( BL35, BLN35, WL81);
sram_cell_6t_3 inst_cell_81_34 ( BL34, BLN34, WL81);
sram_cell_6t_3 inst_cell_81_33 ( BL33, BLN33, WL81);
sram_cell_6t_3 inst_cell_81_32 ( BL32, BLN32, WL81);
sram_cell_6t_3 inst_cell_81_31 ( BL31, BLN31, WL81);
sram_cell_6t_3 inst_cell_81_30 ( BL30, BLN30, WL81);
sram_cell_6t_3 inst_cell_81_29 ( BL29, BLN29, WL81);
sram_cell_6t_3 inst_cell_81_28 ( BL28, BLN28, WL81);
sram_cell_6t_3 inst_cell_81_27 ( BL27, BLN27, WL81);
sram_cell_6t_3 inst_cell_81_26 ( BL26, BLN26, WL81);
sram_cell_6t_3 inst_cell_81_25 ( BL25, BLN25, WL81);
sram_cell_6t_3 inst_cell_81_24 ( BL24, BLN24, WL81);
sram_cell_6t_3 inst_cell_81_23 ( BL23, BLN23, WL81);
sram_cell_6t_3 inst_cell_81_22 ( BL22, BLN22, WL81);
sram_cell_6t_3 inst_cell_81_21 ( BL21, BLN21, WL81);
sram_cell_6t_3 inst_cell_81_20 ( BL20, BLN20, WL81);
sram_cell_6t_3 inst_cell_81_19 ( BL19, BLN19, WL81);
sram_cell_6t_3 inst_cell_81_18 ( BL18, BLN18, WL81);
sram_cell_6t_3 inst_cell_81_17 ( BL17, BLN17, WL81);
sram_cell_6t_3 inst_cell_81_16 ( BL16, BLN16, WL81);
sram_cell_6t_3 inst_cell_81_15 ( BL15, BLN15, WL81);
sram_cell_6t_3 inst_cell_81_14 ( BL14, BLN14, WL81);
sram_cell_6t_3 inst_cell_81_13 ( BL13, BLN13, WL81);
sram_cell_6t_3 inst_cell_81_12 ( BL12, BLN12, WL81);
sram_cell_6t_3 inst_cell_81_11 ( BL11, BLN11, WL81);
sram_cell_6t_3 inst_cell_81_10 ( BL10, BLN10, WL81);
sram_cell_6t_3 inst_cell_81_9 ( BL9, BLN9, WL81);
sram_cell_6t_3 inst_cell_81_8 ( BL8, BLN8, WL81);
sram_cell_6t_3 inst_cell_81_7 ( BL7, BLN7, WL81);
sram_cell_6t_3 inst_cell_81_6 ( BL6, BLN6, WL81);
sram_cell_6t_3 inst_cell_81_5 ( BL5, BLN5, WL81);
sram_cell_6t_3 inst_cell_81_4 ( BL4, BLN4, WL81);
sram_cell_6t_3 inst_cell_81_3 ( BL3, BLN3, WL81);
sram_cell_6t_3 inst_cell_81_2 ( BL2, BLN2, WL81);
sram_cell_6t_3 inst_cell_81_1 ( BL1, BLN1, WL81);
sram_cell_6t_3 inst_cell_81_0 ( BL0, BLN0, WL81);
sram_cell_6t_3 inst_cell_80_127 ( BL127, BLN127, WL80);
sram_cell_6t_3 inst_cell_80_126 ( BL126, BLN126, WL80);
sram_cell_6t_3 inst_cell_80_125 ( BL125, BLN125, WL80);
sram_cell_6t_3 inst_cell_80_124 ( BL124, BLN124, WL80);
sram_cell_6t_3 inst_cell_80_123 ( BL123, BLN123, WL80);
sram_cell_6t_3 inst_cell_80_122 ( BL122, BLN122, WL80);
sram_cell_6t_3 inst_cell_80_121 ( BL121, BLN121, WL80);
sram_cell_6t_3 inst_cell_80_120 ( BL120, BLN120, WL80);
sram_cell_6t_3 inst_cell_80_119 ( BL119, BLN119, WL80);
sram_cell_6t_3 inst_cell_80_118 ( BL118, BLN118, WL80);
sram_cell_6t_3 inst_cell_80_117 ( BL117, BLN117, WL80);
sram_cell_6t_3 inst_cell_80_116 ( BL116, BLN116, WL80);
sram_cell_6t_3 inst_cell_80_115 ( BL115, BLN115, WL80);
sram_cell_6t_3 inst_cell_80_114 ( BL114, BLN114, WL80);
sram_cell_6t_3 inst_cell_80_113 ( BL113, BLN113, WL80);
sram_cell_6t_3 inst_cell_80_112 ( BL112, BLN112, WL80);
sram_cell_6t_3 inst_cell_80_111 ( BL111, BLN111, WL80);
sram_cell_6t_3 inst_cell_80_110 ( BL110, BLN110, WL80);
sram_cell_6t_3 inst_cell_80_109 ( BL109, BLN109, WL80);
sram_cell_6t_3 inst_cell_80_108 ( BL108, BLN108, WL80);
sram_cell_6t_3 inst_cell_80_107 ( BL107, BLN107, WL80);
sram_cell_6t_3 inst_cell_80_106 ( BL106, BLN106, WL80);
sram_cell_6t_3 inst_cell_80_105 ( BL105, BLN105, WL80);
sram_cell_6t_3 inst_cell_80_104 ( BL104, BLN104, WL80);
sram_cell_6t_3 inst_cell_80_103 ( BL103, BLN103, WL80);
sram_cell_6t_3 inst_cell_80_102 ( BL102, BLN102, WL80);
sram_cell_6t_3 inst_cell_80_101 ( BL101, BLN101, WL80);
sram_cell_6t_3 inst_cell_80_100 ( BL100, BLN100, WL80);
sram_cell_6t_3 inst_cell_80_99 ( BL99, BLN99, WL80);
sram_cell_6t_3 inst_cell_80_98 ( BL98, BLN98, WL80);
sram_cell_6t_3 inst_cell_80_97 ( BL97, BLN97, WL80);
sram_cell_6t_3 inst_cell_80_96 ( BL96, BLN96, WL80);
sram_cell_6t_3 inst_cell_80_95 ( BL95, BLN95, WL80);
sram_cell_6t_3 inst_cell_80_94 ( BL94, BLN94, WL80);
sram_cell_6t_3 inst_cell_80_93 ( BL93, BLN93, WL80);
sram_cell_6t_3 inst_cell_80_92 ( BL92, BLN92, WL80);
sram_cell_6t_3 inst_cell_80_91 ( BL91, BLN91, WL80);
sram_cell_6t_3 inst_cell_80_90 ( BL90, BLN90, WL80);
sram_cell_6t_3 inst_cell_80_89 ( BL89, BLN89, WL80);
sram_cell_6t_3 inst_cell_80_88 ( BL88, BLN88, WL80);
sram_cell_6t_3 inst_cell_80_87 ( BL87, BLN87, WL80);
sram_cell_6t_3 inst_cell_80_86 ( BL86, BLN86, WL80);
sram_cell_6t_3 inst_cell_80_85 ( BL85, BLN85, WL80);
sram_cell_6t_3 inst_cell_80_84 ( BL84, BLN84, WL80);
sram_cell_6t_3 inst_cell_80_83 ( BL83, BLN83, WL80);
sram_cell_6t_3 inst_cell_80_82 ( BL82, BLN82, WL80);
sram_cell_6t_3 inst_cell_80_81 ( BL81, BLN81, WL80);
sram_cell_6t_3 inst_cell_80_80 ( BL80, BLN80, WL80);
sram_cell_6t_3 inst_cell_80_79 ( BL79, BLN79, WL80);
sram_cell_6t_3 inst_cell_80_78 ( BL78, BLN78, WL80);
sram_cell_6t_3 inst_cell_80_77 ( BL77, BLN77, WL80);
sram_cell_6t_3 inst_cell_80_76 ( BL76, BLN76, WL80);
sram_cell_6t_3 inst_cell_80_75 ( BL75, BLN75, WL80);
sram_cell_6t_3 inst_cell_80_74 ( BL74, BLN74, WL80);
sram_cell_6t_3 inst_cell_80_73 ( BL73, BLN73, WL80);
sram_cell_6t_3 inst_cell_80_72 ( BL72, BLN72, WL80);
sram_cell_6t_3 inst_cell_80_71 ( BL71, BLN71, WL80);
sram_cell_6t_3 inst_cell_80_70 ( BL70, BLN70, WL80);
sram_cell_6t_3 inst_cell_80_69 ( BL69, BLN69, WL80);
sram_cell_6t_3 inst_cell_80_68 ( BL68, BLN68, WL80);
sram_cell_6t_3 inst_cell_80_67 ( BL67, BLN67, WL80);
sram_cell_6t_3 inst_cell_80_66 ( BL66, BLN66, WL80);
sram_cell_6t_3 inst_cell_80_65 ( BL65, BLN65, WL80);
sram_cell_6t_3 inst_cell_80_64 ( BL64, BLN64, WL80);
sram_cell_6t_3 inst_cell_80_63 ( BL63, BLN63, WL80);
sram_cell_6t_3 inst_cell_80_62 ( BL62, BLN62, WL80);
sram_cell_6t_3 inst_cell_80_61 ( BL61, BLN61, WL80);
sram_cell_6t_3 inst_cell_80_60 ( BL60, BLN60, WL80);
sram_cell_6t_3 inst_cell_80_59 ( BL59, BLN59, WL80);
sram_cell_6t_3 inst_cell_80_58 ( BL58, BLN58, WL80);
sram_cell_6t_3 inst_cell_80_57 ( BL57, BLN57, WL80);
sram_cell_6t_3 inst_cell_80_56 ( BL56, BLN56, WL80);
sram_cell_6t_3 inst_cell_80_55 ( BL55, BLN55, WL80);
sram_cell_6t_3 inst_cell_80_54 ( BL54, BLN54, WL80);
sram_cell_6t_3 inst_cell_80_53 ( BL53, BLN53, WL80);
sram_cell_6t_3 inst_cell_80_52 ( BL52, BLN52, WL80);
sram_cell_6t_3 inst_cell_80_51 ( BL51, BLN51, WL80);
sram_cell_6t_3 inst_cell_80_50 ( BL50, BLN50, WL80);
sram_cell_6t_3 inst_cell_80_49 ( BL49, BLN49, WL80);
sram_cell_6t_3 inst_cell_80_48 ( BL48, BLN48, WL80);
sram_cell_6t_3 inst_cell_80_47 ( BL47, BLN47, WL80);
sram_cell_6t_3 inst_cell_80_46 ( BL46, BLN46, WL80);
sram_cell_6t_3 inst_cell_80_45 ( BL45, BLN45, WL80);
sram_cell_6t_3 inst_cell_80_44 ( BL44, BLN44, WL80);
sram_cell_6t_3 inst_cell_80_43 ( BL43, BLN43, WL80);
sram_cell_6t_3 inst_cell_80_42 ( BL42, BLN42, WL80);
sram_cell_6t_3 inst_cell_80_41 ( BL41, BLN41, WL80);
sram_cell_6t_3 inst_cell_80_40 ( BL40, BLN40, WL80);
sram_cell_6t_3 inst_cell_80_39 ( BL39, BLN39, WL80);
sram_cell_6t_3 inst_cell_80_38 ( BL38, BLN38, WL80);
sram_cell_6t_3 inst_cell_80_37 ( BL37, BLN37, WL80);
sram_cell_6t_3 inst_cell_80_36 ( BL36, BLN36, WL80);
sram_cell_6t_3 inst_cell_80_35 ( BL35, BLN35, WL80);
sram_cell_6t_3 inst_cell_80_34 ( BL34, BLN34, WL80);
sram_cell_6t_3 inst_cell_80_33 ( BL33, BLN33, WL80);
sram_cell_6t_3 inst_cell_80_32 ( BL32, BLN32, WL80);
sram_cell_6t_3 inst_cell_80_31 ( BL31, BLN31, WL80);
sram_cell_6t_3 inst_cell_80_30 ( BL30, BLN30, WL80);
sram_cell_6t_3 inst_cell_80_29 ( BL29, BLN29, WL80);
sram_cell_6t_3 inst_cell_80_28 ( BL28, BLN28, WL80);
sram_cell_6t_3 inst_cell_80_27 ( BL27, BLN27, WL80);
sram_cell_6t_3 inst_cell_80_26 ( BL26, BLN26, WL80);
sram_cell_6t_3 inst_cell_80_25 ( BL25, BLN25, WL80);
sram_cell_6t_3 inst_cell_80_24 ( BL24, BLN24, WL80);
sram_cell_6t_3 inst_cell_80_23 ( BL23, BLN23, WL80);
sram_cell_6t_3 inst_cell_80_22 ( BL22, BLN22, WL80);
sram_cell_6t_3 inst_cell_80_21 ( BL21, BLN21, WL80);
sram_cell_6t_3 inst_cell_80_20 ( BL20, BLN20, WL80);
sram_cell_6t_3 inst_cell_80_19 ( BL19, BLN19, WL80);
sram_cell_6t_3 inst_cell_80_18 ( BL18, BLN18, WL80);
sram_cell_6t_3 inst_cell_80_17 ( BL17, BLN17, WL80);
sram_cell_6t_3 inst_cell_80_16 ( BL16, BLN16, WL80);
sram_cell_6t_3 inst_cell_80_15 ( BL15, BLN15, WL80);
sram_cell_6t_3 inst_cell_80_14 ( BL14, BLN14, WL80);
sram_cell_6t_3 inst_cell_80_13 ( BL13, BLN13, WL80);
sram_cell_6t_3 inst_cell_80_12 ( BL12, BLN12, WL80);
sram_cell_6t_3 inst_cell_80_11 ( BL11, BLN11, WL80);
sram_cell_6t_3 inst_cell_80_10 ( BL10, BLN10, WL80);
sram_cell_6t_3 inst_cell_80_9 ( BL9, BLN9, WL80);
sram_cell_6t_3 inst_cell_80_8 ( BL8, BLN8, WL80);
sram_cell_6t_3 inst_cell_80_7 ( BL7, BLN7, WL80);
sram_cell_6t_3 inst_cell_80_6 ( BL6, BLN6, WL80);
sram_cell_6t_3 inst_cell_80_5 ( BL5, BLN5, WL80);
sram_cell_6t_3 inst_cell_80_4 ( BL4, BLN4, WL80);
sram_cell_6t_3 inst_cell_80_3 ( BL3, BLN3, WL80);
sram_cell_6t_3 inst_cell_80_2 ( BL2, BLN2, WL80);
sram_cell_6t_3 inst_cell_80_1 ( BL1, BLN1, WL80);
sram_cell_6t_3 inst_cell_80_0 ( BL0, BLN0, WL80);
sram_cell_6t_3 inst_cell_79_127 ( BL127, BLN127, WL79);
sram_cell_6t_3 inst_cell_79_126 ( BL126, BLN126, WL79);
sram_cell_6t_3 inst_cell_79_125 ( BL125, BLN125, WL79);
sram_cell_6t_3 inst_cell_79_124 ( BL124, BLN124, WL79);
sram_cell_6t_3 inst_cell_79_123 ( BL123, BLN123, WL79);
sram_cell_6t_3 inst_cell_79_122 ( BL122, BLN122, WL79);
sram_cell_6t_3 inst_cell_79_121 ( BL121, BLN121, WL79);
sram_cell_6t_3 inst_cell_79_120 ( BL120, BLN120, WL79);
sram_cell_6t_3 inst_cell_79_119 ( BL119, BLN119, WL79);
sram_cell_6t_3 inst_cell_79_118 ( BL118, BLN118, WL79);
sram_cell_6t_3 inst_cell_79_117 ( BL117, BLN117, WL79);
sram_cell_6t_3 inst_cell_79_116 ( BL116, BLN116, WL79);
sram_cell_6t_3 inst_cell_79_115 ( BL115, BLN115, WL79);
sram_cell_6t_3 inst_cell_79_114 ( BL114, BLN114, WL79);
sram_cell_6t_3 inst_cell_79_113 ( BL113, BLN113, WL79);
sram_cell_6t_3 inst_cell_79_112 ( BL112, BLN112, WL79);
sram_cell_6t_3 inst_cell_79_111 ( BL111, BLN111, WL79);
sram_cell_6t_3 inst_cell_79_110 ( BL110, BLN110, WL79);
sram_cell_6t_3 inst_cell_79_109 ( BL109, BLN109, WL79);
sram_cell_6t_3 inst_cell_79_108 ( BL108, BLN108, WL79);
sram_cell_6t_3 inst_cell_79_107 ( BL107, BLN107, WL79);
sram_cell_6t_3 inst_cell_79_106 ( BL106, BLN106, WL79);
sram_cell_6t_3 inst_cell_79_105 ( BL105, BLN105, WL79);
sram_cell_6t_3 inst_cell_79_104 ( BL104, BLN104, WL79);
sram_cell_6t_3 inst_cell_79_103 ( BL103, BLN103, WL79);
sram_cell_6t_3 inst_cell_79_102 ( BL102, BLN102, WL79);
sram_cell_6t_3 inst_cell_79_101 ( BL101, BLN101, WL79);
sram_cell_6t_3 inst_cell_79_100 ( BL100, BLN100, WL79);
sram_cell_6t_3 inst_cell_79_99 ( BL99, BLN99, WL79);
sram_cell_6t_3 inst_cell_79_98 ( BL98, BLN98, WL79);
sram_cell_6t_3 inst_cell_79_97 ( BL97, BLN97, WL79);
sram_cell_6t_3 inst_cell_79_96 ( BL96, BLN96, WL79);
sram_cell_6t_3 inst_cell_79_95 ( BL95, BLN95, WL79);
sram_cell_6t_3 inst_cell_79_94 ( BL94, BLN94, WL79);
sram_cell_6t_3 inst_cell_79_93 ( BL93, BLN93, WL79);
sram_cell_6t_3 inst_cell_79_92 ( BL92, BLN92, WL79);
sram_cell_6t_3 inst_cell_79_91 ( BL91, BLN91, WL79);
sram_cell_6t_3 inst_cell_79_90 ( BL90, BLN90, WL79);
sram_cell_6t_3 inst_cell_79_89 ( BL89, BLN89, WL79);
sram_cell_6t_3 inst_cell_79_88 ( BL88, BLN88, WL79);
sram_cell_6t_3 inst_cell_79_87 ( BL87, BLN87, WL79);
sram_cell_6t_3 inst_cell_79_86 ( BL86, BLN86, WL79);
sram_cell_6t_3 inst_cell_79_85 ( BL85, BLN85, WL79);
sram_cell_6t_3 inst_cell_79_84 ( BL84, BLN84, WL79);
sram_cell_6t_3 inst_cell_79_83 ( BL83, BLN83, WL79);
sram_cell_6t_3 inst_cell_79_82 ( BL82, BLN82, WL79);
sram_cell_6t_3 inst_cell_79_81 ( BL81, BLN81, WL79);
sram_cell_6t_3 inst_cell_79_80 ( BL80, BLN80, WL79);
sram_cell_6t_3 inst_cell_79_79 ( BL79, BLN79, WL79);
sram_cell_6t_3 inst_cell_79_78 ( BL78, BLN78, WL79);
sram_cell_6t_3 inst_cell_79_77 ( BL77, BLN77, WL79);
sram_cell_6t_3 inst_cell_79_76 ( BL76, BLN76, WL79);
sram_cell_6t_3 inst_cell_79_75 ( BL75, BLN75, WL79);
sram_cell_6t_3 inst_cell_79_74 ( BL74, BLN74, WL79);
sram_cell_6t_3 inst_cell_79_73 ( BL73, BLN73, WL79);
sram_cell_6t_3 inst_cell_79_72 ( BL72, BLN72, WL79);
sram_cell_6t_3 inst_cell_79_71 ( BL71, BLN71, WL79);
sram_cell_6t_3 inst_cell_79_70 ( BL70, BLN70, WL79);
sram_cell_6t_3 inst_cell_79_69 ( BL69, BLN69, WL79);
sram_cell_6t_3 inst_cell_79_68 ( BL68, BLN68, WL79);
sram_cell_6t_3 inst_cell_79_67 ( BL67, BLN67, WL79);
sram_cell_6t_3 inst_cell_79_66 ( BL66, BLN66, WL79);
sram_cell_6t_3 inst_cell_79_65 ( BL65, BLN65, WL79);
sram_cell_6t_3 inst_cell_79_64 ( BL64, BLN64, WL79);
sram_cell_6t_3 inst_cell_79_63 ( BL63, BLN63, WL79);
sram_cell_6t_3 inst_cell_79_62 ( BL62, BLN62, WL79);
sram_cell_6t_3 inst_cell_79_61 ( BL61, BLN61, WL79);
sram_cell_6t_3 inst_cell_79_60 ( BL60, BLN60, WL79);
sram_cell_6t_3 inst_cell_79_59 ( BL59, BLN59, WL79);
sram_cell_6t_3 inst_cell_79_58 ( BL58, BLN58, WL79);
sram_cell_6t_3 inst_cell_79_57 ( BL57, BLN57, WL79);
sram_cell_6t_3 inst_cell_79_56 ( BL56, BLN56, WL79);
sram_cell_6t_3 inst_cell_79_55 ( BL55, BLN55, WL79);
sram_cell_6t_3 inst_cell_79_54 ( BL54, BLN54, WL79);
sram_cell_6t_3 inst_cell_79_53 ( BL53, BLN53, WL79);
sram_cell_6t_3 inst_cell_79_52 ( BL52, BLN52, WL79);
sram_cell_6t_3 inst_cell_79_51 ( BL51, BLN51, WL79);
sram_cell_6t_3 inst_cell_79_50 ( BL50, BLN50, WL79);
sram_cell_6t_3 inst_cell_79_49 ( BL49, BLN49, WL79);
sram_cell_6t_3 inst_cell_79_48 ( BL48, BLN48, WL79);
sram_cell_6t_3 inst_cell_79_47 ( BL47, BLN47, WL79);
sram_cell_6t_3 inst_cell_79_46 ( BL46, BLN46, WL79);
sram_cell_6t_3 inst_cell_79_45 ( BL45, BLN45, WL79);
sram_cell_6t_3 inst_cell_79_44 ( BL44, BLN44, WL79);
sram_cell_6t_3 inst_cell_79_43 ( BL43, BLN43, WL79);
sram_cell_6t_3 inst_cell_79_42 ( BL42, BLN42, WL79);
sram_cell_6t_3 inst_cell_79_41 ( BL41, BLN41, WL79);
sram_cell_6t_3 inst_cell_79_40 ( BL40, BLN40, WL79);
sram_cell_6t_3 inst_cell_79_39 ( BL39, BLN39, WL79);
sram_cell_6t_3 inst_cell_79_38 ( BL38, BLN38, WL79);
sram_cell_6t_3 inst_cell_79_37 ( BL37, BLN37, WL79);
sram_cell_6t_3 inst_cell_79_36 ( BL36, BLN36, WL79);
sram_cell_6t_3 inst_cell_79_35 ( BL35, BLN35, WL79);
sram_cell_6t_3 inst_cell_79_34 ( BL34, BLN34, WL79);
sram_cell_6t_3 inst_cell_79_33 ( BL33, BLN33, WL79);
sram_cell_6t_3 inst_cell_79_32 ( BL32, BLN32, WL79);
sram_cell_6t_3 inst_cell_79_31 ( BL31, BLN31, WL79);
sram_cell_6t_3 inst_cell_79_30 ( BL30, BLN30, WL79);
sram_cell_6t_3 inst_cell_79_29 ( BL29, BLN29, WL79);
sram_cell_6t_3 inst_cell_79_28 ( BL28, BLN28, WL79);
sram_cell_6t_3 inst_cell_79_27 ( BL27, BLN27, WL79);
sram_cell_6t_3 inst_cell_79_26 ( BL26, BLN26, WL79);
sram_cell_6t_3 inst_cell_79_25 ( BL25, BLN25, WL79);
sram_cell_6t_3 inst_cell_79_24 ( BL24, BLN24, WL79);
sram_cell_6t_3 inst_cell_79_23 ( BL23, BLN23, WL79);
sram_cell_6t_3 inst_cell_79_22 ( BL22, BLN22, WL79);
sram_cell_6t_3 inst_cell_79_21 ( BL21, BLN21, WL79);
sram_cell_6t_3 inst_cell_79_20 ( BL20, BLN20, WL79);
sram_cell_6t_3 inst_cell_79_19 ( BL19, BLN19, WL79);
sram_cell_6t_3 inst_cell_79_18 ( BL18, BLN18, WL79);
sram_cell_6t_3 inst_cell_79_17 ( BL17, BLN17, WL79);
sram_cell_6t_3 inst_cell_79_16 ( BL16, BLN16, WL79);
sram_cell_6t_3 inst_cell_79_15 ( BL15, BLN15, WL79);
sram_cell_6t_3 inst_cell_79_14 ( BL14, BLN14, WL79);
sram_cell_6t_3 inst_cell_79_13 ( BL13, BLN13, WL79);
sram_cell_6t_3 inst_cell_79_12 ( BL12, BLN12, WL79);
sram_cell_6t_3 inst_cell_79_11 ( BL11, BLN11, WL79);
sram_cell_6t_3 inst_cell_79_10 ( BL10, BLN10, WL79);
sram_cell_6t_3 inst_cell_79_9 ( BL9, BLN9, WL79);
sram_cell_6t_3 inst_cell_79_8 ( BL8, BLN8, WL79);
sram_cell_6t_3 inst_cell_79_7 ( BL7, BLN7, WL79);
sram_cell_6t_3 inst_cell_79_6 ( BL6, BLN6, WL79);
sram_cell_6t_3 inst_cell_79_5 ( BL5, BLN5, WL79);
sram_cell_6t_3 inst_cell_79_4 ( BL4, BLN4, WL79);
sram_cell_6t_3 inst_cell_79_3 ( BL3, BLN3, WL79);
sram_cell_6t_3 inst_cell_79_2 ( BL2, BLN2, WL79);
sram_cell_6t_3 inst_cell_79_1 ( BL1, BLN1, WL79);
sram_cell_6t_3 inst_cell_79_0 ( BL0, BLN0, WL79);
sram_cell_6t_3 inst_cell_78_127 ( BL127, BLN127, WL78);
sram_cell_6t_3 inst_cell_78_126 ( BL126, BLN126, WL78);
sram_cell_6t_3 inst_cell_78_125 ( BL125, BLN125, WL78);
sram_cell_6t_3 inst_cell_78_124 ( BL124, BLN124, WL78);
sram_cell_6t_3 inst_cell_78_123 ( BL123, BLN123, WL78);
sram_cell_6t_3 inst_cell_78_122 ( BL122, BLN122, WL78);
sram_cell_6t_3 inst_cell_78_121 ( BL121, BLN121, WL78);
sram_cell_6t_3 inst_cell_78_120 ( BL120, BLN120, WL78);
sram_cell_6t_3 inst_cell_78_119 ( BL119, BLN119, WL78);
sram_cell_6t_3 inst_cell_78_118 ( BL118, BLN118, WL78);
sram_cell_6t_3 inst_cell_78_117 ( BL117, BLN117, WL78);
sram_cell_6t_3 inst_cell_78_116 ( BL116, BLN116, WL78);
sram_cell_6t_3 inst_cell_78_115 ( BL115, BLN115, WL78);
sram_cell_6t_3 inst_cell_78_114 ( BL114, BLN114, WL78);
sram_cell_6t_3 inst_cell_78_113 ( BL113, BLN113, WL78);
sram_cell_6t_3 inst_cell_78_112 ( BL112, BLN112, WL78);
sram_cell_6t_3 inst_cell_78_111 ( BL111, BLN111, WL78);
sram_cell_6t_3 inst_cell_78_110 ( BL110, BLN110, WL78);
sram_cell_6t_3 inst_cell_78_109 ( BL109, BLN109, WL78);
sram_cell_6t_3 inst_cell_78_108 ( BL108, BLN108, WL78);
sram_cell_6t_3 inst_cell_78_107 ( BL107, BLN107, WL78);
sram_cell_6t_3 inst_cell_78_106 ( BL106, BLN106, WL78);
sram_cell_6t_3 inst_cell_78_105 ( BL105, BLN105, WL78);
sram_cell_6t_3 inst_cell_78_104 ( BL104, BLN104, WL78);
sram_cell_6t_3 inst_cell_78_103 ( BL103, BLN103, WL78);
sram_cell_6t_3 inst_cell_78_102 ( BL102, BLN102, WL78);
sram_cell_6t_3 inst_cell_78_101 ( BL101, BLN101, WL78);
sram_cell_6t_3 inst_cell_78_100 ( BL100, BLN100, WL78);
sram_cell_6t_3 inst_cell_78_99 ( BL99, BLN99, WL78);
sram_cell_6t_3 inst_cell_78_98 ( BL98, BLN98, WL78);
sram_cell_6t_3 inst_cell_78_97 ( BL97, BLN97, WL78);
sram_cell_6t_3 inst_cell_78_96 ( BL96, BLN96, WL78);
sram_cell_6t_3 inst_cell_78_95 ( BL95, BLN95, WL78);
sram_cell_6t_3 inst_cell_78_94 ( BL94, BLN94, WL78);
sram_cell_6t_3 inst_cell_78_93 ( BL93, BLN93, WL78);
sram_cell_6t_3 inst_cell_78_92 ( BL92, BLN92, WL78);
sram_cell_6t_3 inst_cell_78_91 ( BL91, BLN91, WL78);
sram_cell_6t_3 inst_cell_78_90 ( BL90, BLN90, WL78);
sram_cell_6t_3 inst_cell_78_89 ( BL89, BLN89, WL78);
sram_cell_6t_3 inst_cell_78_88 ( BL88, BLN88, WL78);
sram_cell_6t_3 inst_cell_78_87 ( BL87, BLN87, WL78);
sram_cell_6t_3 inst_cell_78_86 ( BL86, BLN86, WL78);
sram_cell_6t_3 inst_cell_78_85 ( BL85, BLN85, WL78);
sram_cell_6t_3 inst_cell_78_84 ( BL84, BLN84, WL78);
sram_cell_6t_3 inst_cell_78_83 ( BL83, BLN83, WL78);
sram_cell_6t_3 inst_cell_78_82 ( BL82, BLN82, WL78);
sram_cell_6t_3 inst_cell_78_81 ( BL81, BLN81, WL78);
sram_cell_6t_3 inst_cell_78_80 ( BL80, BLN80, WL78);
sram_cell_6t_3 inst_cell_78_79 ( BL79, BLN79, WL78);
sram_cell_6t_3 inst_cell_78_78 ( BL78, BLN78, WL78);
sram_cell_6t_3 inst_cell_78_77 ( BL77, BLN77, WL78);
sram_cell_6t_3 inst_cell_78_76 ( BL76, BLN76, WL78);
sram_cell_6t_3 inst_cell_78_75 ( BL75, BLN75, WL78);
sram_cell_6t_3 inst_cell_78_74 ( BL74, BLN74, WL78);
sram_cell_6t_3 inst_cell_78_73 ( BL73, BLN73, WL78);
sram_cell_6t_3 inst_cell_78_72 ( BL72, BLN72, WL78);
sram_cell_6t_3 inst_cell_78_71 ( BL71, BLN71, WL78);
sram_cell_6t_3 inst_cell_78_70 ( BL70, BLN70, WL78);
sram_cell_6t_3 inst_cell_78_69 ( BL69, BLN69, WL78);
sram_cell_6t_3 inst_cell_78_68 ( BL68, BLN68, WL78);
sram_cell_6t_3 inst_cell_78_67 ( BL67, BLN67, WL78);
sram_cell_6t_3 inst_cell_78_66 ( BL66, BLN66, WL78);
sram_cell_6t_3 inst_cell_78_65 ( BL65, BLN65, WL78);
sram_cell_6t_3 inst_cell_78_64 ( BL64, BLN64, WL78);
sram_cell_6t_3 inst_cell_78_63 ( BL63, BLN63, WL78);
sram_cell_6t_3 inst_cell_78_62 ( BL62, BLN62, WL78);
sram_cell_6t_3 inst_cell_78_61 ( BL61, BLN61, WL78);
sram_cell_6t_3 inst_cell_78_60 ( BL60, BLN60, WL78);
sram_cell_6t_3 inst_cell_78_59 ( BL59, BLN59, WL78);
sram_cell_6t_3 inst_cell_78_58 ( BL58, BLN58, WL78);
sram_cell_6t_3 inst_cell_78_57 ( BL57, BLN57, WL78);
sram_cell_6t_3 inst_cell_78_56 ( BL56, BLN56, WL78);
sram_cell_6t_3 inst_cell_78_55 ( BL55, BLN55, WL78);
sram_cell_6t_3 inst_cell_78_54 ( BL54, BLN54, WL78);
sram_cell_6t_3 inst_cell_78_53 ( BL53, BLN53, WL78);
sram_cell_6t_3 inst_cell_78_52 ( BL52, BLN52, WL78);
sram_cell_6t_3 inst_cell_78_51 ( BL51, BLN51, WL78);
sram_cell_6t_3 inst_cell_78_50 ( BL50, BLN50, WL78);
sram_cell_6t_3 inst_cell_78_49 ( BL49, BLN49, WL78);
sram_cell_6t_3 inst_cell_78_48 ( BL48, BLN48, WL78);
sram_cell_6t_3 inst_cell_78_47 ( BL47, BLN47, WL78);
sram_cell_6t_3 inst_cell_78_46 ( BL46, BLN46, WL78);
sram_cell_6t_3 inst_cell_78_45 ( BL45, BLN45, WL78);
sram_cell_6t_3 inst_cell_78_44 ( BL44, BLN44, WL78);
sram_cell_6t_3 inst_cell_78_43 ( BL43, BLN43, WL78);
sram_cell_6t_3 inst_cell_78_42 ( BL42, BLN42, WL78);
sram_cell_6t_3 inst_cell_78_41 ( BL41, BLN41, WL78);
sram_cell_6t_3 inst_cell_78_40 ( BL40, BLN40, WL78);
sram_cell_6t_3 inst_cell_78_39 ( BL39, BLN39, WL78);
sram_cell_6t_3 inst_cell_78_38 ( BL38, BLN38, WL78);
sram_cell_6t_3 inst_cell_78_37 ( BL37, BLN37, WL78);
sram_cell_6t_3 inst_cell_78_36 ( BL36, BLN36, WL78);
sram_cell_6t_3 inst_cell_78_35 ( BL35, BLN35, WL78);
sram_cell_6t_3 inst_cell_78_34 ( BL34, BLN34, WL78);
sram_cell_6t_3 inst_cell_78_33 ( BL33, BLN33, WL78);
sram_cell_6t_3 inst_cell_78_32 ( BL32, BLN32, WL78);
sram_cell_6t_3 inst_cell_78_31 ( BL31, BLN31, WL78);
sram_cell_6t_3 inst_cell_78_30 ( BL30, BLN30, WL78);
sram_cell_6t_3 inst_cell_78_29 ( BL29, BLN29, WL78);
sram_cell_6t_3 inst_cell_78_28 ( BL28, BLN28, WL78);
sram_cell_6t_3 inst_cell_78_27 ( BL27, BLN27, WL78);
sram_cell_6t_3 inst_cell_78_26 ( BL26, BLN26, WL78);
sram_cell_6t_3 inst_cell_78_25 ( BL25, BLN25, WL78);
sram_cell_6t_3 inst_cell_78_24 ( BL24, BLN24, WL78);
sram_cell_6t_3 inst_cell_78_23 ( BL23, BLN23, WL78);
sram_cell_6t_3 inst_cell_78_22 ( BL22, BLN22, WL78);
sram_cell_6t_3 inst_cell_78_21 ( BL21, BLN21, WL78);
sram_cell_6t_3 inst_cell_78_20 ( BL20, BLN20, WL78);
sram_cell_6t_3 inst_cell_78_19 ( BL19, BLN19, WL78);
sram_cell_6t_3 inst_cell_78_18 ( BL18, BLN18, WL78);
sram_cell_6t_3 inst_cell_78_17 ( BL17, BLN17, WL78);
sram_cell_6t_3 inst_cell_78_16 ( BL16, BLN16, WL78);
sram_cell_6t_3 inst_cell_78_15 ( BL15, BLN15, WL78);
sram_cell_6t_3 inst_cell_78_14 ( BL14, BLN14, WL78);
sram_cell_6t_3 inst_cell_78_13 ( BL13, BLN13, WL78);
sram_cell_6t_3 inst_cell_78_12 ( BL12, BLN12, WL78);
sram_cell_6t_3 inst_cell_78_11 ( BL11, BLN11, WL78);
sram_cell_6t_3 inst_cell_78_10 ( BL10, BLN10, WL78);
sram_cell_6t_3 inst_cell_78_9 ( BL9, BLN9, WL78);
sram_cell_6t_3 inst_cell_78_8 ( BL8, BLN8, WL78);
sram_cell_6t_3 inst_cell_78_7 ( BL7, BLN7, WL78);
sram_cell_6t_3 inst_cell_78_6 ( BL6, BLN6, WL78);
sram_cell_6t_3 inst_cell_78_5 ( BL5, BLN5, WL78);
sram_cell_6t_3 inst_cell_78_4 ( BL4, BLN4, WL78);
sram_cell_6t_3 inst_cell_78_3 ( BL3, BLN3, WL78);
sram_cell_6t_3 inst_cell_78_2 ( BL2, BLN2, WL78);
sram_cell_6t_3 inst_cell_78_1 ( BL1, BLN1, WL78);
sram_cell_6t_3 inst_cell_78_0 ( BL0, BLN0, WL78);
sram_cell_6t_3 inst_cell_77_127 ( BL127, BLN127, WL77);
sram_cell_6t_3 inst_cell_77_126 ( BL126, BLN126, WL77);
sram_cell_6t_3 inst_cell_77_125 ( BL125, BLN125, WL77);
sram_cell_6t_3 inst_cell_77_124 ( BL124, BLN124, WL77);
sram_cell_6t_3 inst_cell_77_123 ( BL123, BLN123, WL77);
sram_cell_6t_3 inst_cell_77_122 ( BL122, BLN122, WL77);
sram_cell_6t_3 inst_cell_77_121 ( BL121, BLN121, WL77);
sram_cell_6t_3 inst_cell_77_120 ( BL120, BLN120, WL77);
sram_cell_6t_3 inst_cell_77_119 ( BL119, BLN119, WL77);
sram_cell_6t_3 inst_cell_77_118 ( BL118, BLN118, WL77);
sram_cell_6t_3 inst_cell_77_117 ( BL117, BLN117, WL77);
sram_cell_6t_3 inst_cell_77_116 ( BL116, BLN116, WL77);
sram_cell_6t_3 inst_cell_77_115 ( BL115, BLN115, WL77);
sram_cell_6t_3 inst_cell_77_114 ( BL114, BLN114, WL77);
sram_cell_6t_3 inst_cell_77_113 ( BL113, BLN113, WL77);
sram_cell_6t_3 inst_cell_77_112 ( BL112, BLN112, WL77);
sram_cell_6t_3 inst_cell_77_111 ( BL111, BLN111, WL77);
sram_cell_6t_3 inst_cell_77_110 ( BL110, BLN110, WL77);
sram_cell_6t_3 inst_cell_77_109 ( BL109, BLN109, WL77);
sram_cell_6t_3 inst_cell_77_108 ( BL108, BLN108, WL77);
sram_cell_6t_3 inst_cell_77_107 ( BL107, BLN107, WL77);
sram_cell_6t_3 inst_cell_77_106 ( BL106, BLN106, WL77);
sram_cell_6t_3 inst_cell_77_105 ( BL105, BLN105, WL77);
sram_cell_6t_3 inst_cell_77_104 ( BL104, BLN104, WL77);
sram_cell_6t_3 inst_cell_77_103 ( BL103, BLN103, WL77);
sram_cell_6t_3 inst_cell_77_102 ( BL102, BLN102, WL77);
sram_cell_6t_3 inst_cell_77_101 ( BL101, BLN101, WL77);
sram_cell_6t_3 inst_cell_77_100 ( BL100, BLN100, WL77);
sram_cell_6t_3 inst_cell_77_99 ( BL99, BLN99, WL77);
sram_cell_6t_3 inst_cell_77_98 ( BL98, BLN98, WL77);
sram_cell_6t_3 inst_cell_77_97 ( BL97, BLN97, WL77);
sram_cell_6t_3 inst_cell_77_96 ( BL96, BLN96, WL77);
sram_cell_6t_3 inst_cell_77_95 ( BL95, BLN95, WL77);
sram_cell_6t_3 inst_cell_77_94 ( BL94, BLN94, WL77);
sram_cell_6t_3 inst_cell_77_93 ( BL93, BLN93, WL77);
sram_cell_6t_3 inst_cell_77_92 ( BL92, BLN92, WL77);
sram_cell_6t_3 inst_cell_77_91 ( BL91, BLN91, WL77);
sram_cell_6t_3 inst_cell_77_90 ( BL90, BLN90, WL77);
sram_cell_6t_3 inst_cell_77_89 ( BL89, BLN89, WL77);
sram_cell_6t_3 inst_cell_77_88 ( BL88, BLN88, WL77);
sram_cell_6t_3 inst_cell_77_87 ( BL87, BLN87, WL77);
sram_cell_6t_3 inst_cell_77_86 ( BL86, BLN86, WL77);
sram_cell_6t_3 inst_cell_77_85 ( BL85, BLN85, WL77);
sram_cell_6t_3 inst_cell_77_84 ( BL84, BLN84, WL77);
sram_cell_6t_3 inst_cell_77_83 ( BL83, BLN83, WL77);
sram_cell_6t_3 inst_cell_77_82 ( BL82, BLN82, WL77);
sram_cell_6t_3 inst_cell_77_81 ( BL81, BLN81, WL77);
sram_cell_6t_3 inst_cell_77_80 ( BL80, BLN80, WL77);
sram_cell_6t_3 inst_cell_77_79 ( BL79, BLN79, WL77);
sram_cell_6t_3 inst_cell_77_78 ( BL78, BLN78, WL77);
sram_cell_6t_3 inst_cell_77_77 ( BL77, BLN77, WL77);
sram_cell_6t_3 inst_cell_77_76 ( BL76, BLN76, WL77);
sram_cell_6t_3 inst_cell_77_75 ( BL75, BLN75, WL77);
sram_cell_6t_3 inst_cell_77_74 ( BL74, BLN74, WL77);
sram_cell_6t_3 inst_cell_77_73 ( BL73, BLN73, WL77);
sram_cell_6t_3 inst_cell_77_72 ( BL72, BLN72, WL77);
sram_cell_6t_3 inst_cell_77_71 ( BL71, BLN71, WL77);
sram_cell_6t_3 inst_cell_77_70 ( BL70, BLN70, WL77);
sram_cell_6t_3 inst_cell_77_69 ( BL69, BLN69, WL77);
sram_cell_6t_3 inst_cell_77_68 ( BL68, BLN68, WL77);
sram_cell_6t_3 inst_cell_77_67 ( BL67, BLN67, WL77);
sram_cell_6t_3 inst_cell_77_66 ( BL66, BLN66, WL77);
sram_cell_6t_3 inst_cell_77_65 ( BL65, BLN65, WL77);
sram_cell_6t_3 inst_cell_77_64 ( BL64, BLN64, WL77);
sram_cell_6t_3 inst_cell_77_63 ( BL63, BLN63, WL77);
sram_cell_6t_3 inst_cell_77_62 ( BL62, BLN62, WL77);
sram_cell_6t_3 inst_cell_77_61 ( BL61, BLN61, WL77);
sram_cell_6t_3 inst_cell_77_60 ( BL60, BLN60, WL77);
sram_cell_6t_3 inst_cell_77_59 ( BL59, BLN59, WL77);
sram_cell_6t_3 inst_cell_77_58 ( BL58, BLN58, WL77);
sram_cell_6t_3 inst_cell_77_57 ( BL57, BLN57, WL77);
sram_cell_6t_3 inst_cell_77_56 ( BL56, BLN56, WL77);
sram_cell_6t_3 inst_cell_77_55 ( BL55, BLN55, WL77);
sram_cell_6t_3 inst_cell_77_54 ( BL54, BLN54, WL77);
sram_cell_6t_3 inst_cell_77_53 ( BL53, BLN53, WL77);
sram_cell_6t_3 inst_cell_77_52 ( BL52, BLN52, WL77);
sram_cell_6t_3 inst_cell_77_51 ( BL51, BLN51, WL77);
sram_cell_6t_3 inst_cell_77_50 ( BL50, BLN50, WL77);
sram_cell_6t_3 inst_cell_77_49 ( BL49, BLN49, WL77);
sram_cell_6t_3 inst_cell_77_48 ( BL48, BLN48, WL77);
sram_cell_6t_3 inst_cell_77_47 ( BL47, BLN47, WL77);
sram_cell_6t_3 inst_cell_77_46 ( BL46, BLN46, WL77);
sram_cell_6t_3 inst_cell_77_45 ( BL45, BLN45, WL77);
sram_cell_6t_3 inst_cell_77_44 ( BL44, BLN44, WL77);
sram_cell_6t_3 inst_cell_77_43 ( BL43, BLN43, WL77);
sram_cell_6t_3 inst_cell_77_42 ( BL42, BLN42, WL77);
sram_cell_6t_3 inst_cell_77_41 ( BL41, BLN41, WL77);
sram_cell_6t_3 inst_cell_77_40 ( BL40, BLN40, WL77);
sram_cell_6t_3 inst_cell_77_39 ( BL39, BLN39, WL77);
sram_cell_6t_3 inst_cell_77_38 ( BL38, BLN38, WL77);
sram_cell_6t_3 inst_cell_77_37 ( BL37, BLN37, WL77);
sram_cell_6t_3 inst_cell_77_36 ( BL36, BLN36, WL77);
sram_cell_6t_3 inst_cell_77_35 ( BL35, BLN35, WL77);
sram_cell_6t_3 inst_cell_77_34 ( BL34, BLN34, WL77);
sram_cell_6t_3 inst_cell_77_33 ( BL33, BLN33, WL77);
sram_cell_6t_3 inst_cell_77_32 ( BL32, BLN32, WL77);
sram_cell_6t_3 inst_cell_77_31 ( BL31, BLN31, WL77);
sram_cell_6t_3 inst_cell_77_30 ( BL30, BLN30, WL77);
sram_cell_6t_3 inst_cell_77_29 ( BL29, BLN29, WL77);
sram_cell_6t_3 inst_cell_77_28 ( BL28, BLN28, WL77);
sram_cell_6t_3 inst_cell_77_27 ( BL27, BLN27, WL77);
sram_cell_6t_3 inst_cell_77_26 ( BL26, BLN26, WL77);
sram_cell_6t_3 inst_cell_77_25 ( BL25, BLN25, WL77);
sram_cell_6t_3 inst_cell_77_24 ( BL24, BLN24, WL77);
sram_cell_6t_3 inst_cell_77_23 ( BL23, BLN23, WL77);
sram_cell_6t_3 inst_cell_77_22 ( BL22, BLN22, WL77);
sram_cell_6t_3 inst_cell_77_21 ( BL21, BLN21, WL77);
sram_cell_6t_3 inst_cell_77_20 ( BL20, BLN20, WL77);
sram_cell_6t_3 inst_cell_77_19 ( BL19, BLN19, WL77);
sram_cell_6t_3 inst_cell_77_18 ( BL18, BLN18, WL77);
sram_cell_6t_3 inst_cell_77_17 ( BL17, BLN17, WL77);
sram_cell_6t_3 inst_cell_77_16 ( BL16, BLN16, WL77);
sram_cell_6t_3 inst_cell_77_15 ( BL15, BLN15, WL77);
sram_cell_6t_3 inst_cell_77_14 ( BL14, BLN14, WL77);
sram_cell_6t_3 inst_cell_77_13 ( BL13, BLN13, WL77);
sram_cell_6t_3 inst_cell_77_12 ( BL12, BLN12, WL77);
sram_cell_6t_3 inst_cell_77_11 ( BL11, BLN11, WL77);
sram_cell_6t_3 inst_cell_77_10 ( BL10, BLN10, WL77);
sram_cell_6t_3 inst_cell_77_9 ( BL9, BLN9, WL77);
sram_cell_6t_3 inst_cell_77_8 ( BL8, BLN8, WL77);
sram_cell_6t_3 inst_cell_77_7 ( BL7, BLN7, WL77);
sram_cell_6t_3 inst_cell_77_6 ( BL6, BLN6, WL77);
sram_cell_6t_3 inst_cell_77_5 ( BL5, BLN5, WL77);
sram_cell_6t_3 inst_cell_77_4 ( BL4, BLN4, WL77);
sram_cell_6t_3 inst_cell_77_3 ( BL3, BLN3, WL77);
sram_cell_6t_3 inst_cell_77_2 ( BL2, BLN2, WL77);
sram_cell_6t_3 inst_cell_77_1 ( BL1, BLN1, WL77);
sram_cell_6t_3 inst_cell_77_0 ( BL0, BLN0, WL77);
sram_cell_6t_3 inst_cell_76_127 ( BL127, BLN127, WL76);
sram_cell_6t_3 inst_cell_76_126 ( BL126, BLN126, WL76);
sram_cell_6t_3 inst_cell_76_125 ( BL125, BLN125, WL76);
sram_cell_6t_3 inst_cell_76_124 ( BL124, BLN124, WL76);
sram_cell_6t_3 inst_cell_76_123 ( BL123, BLN123, WL76);
sram_cell_6t_3 inst_cell_76_122 ( BL122, BLN122, WL76);
sram_cell_6t_3 inst_cell_76_121 ( BL121, BLN121, WL76);
sram_cell_6t_3 inst_cell_76_120 ( BL120, BLN120, WL76);
sram_cell_6t_3 inst_cell_76_119 ( BL119, BLN119, WL76);
sram_cell_6t_3 inst_cell_76_118 ( BL118, BLN118, WL76);
sram_cell_6t_3 inst_cell_76_117 ( BL117, BLN117, WL76);
sram_cell_6t_3 inst_cell_76_116 ( BL116, BLN116, WL76);
sram_cell_6t_3 inst_cell_76_115 ( BL115, BLN115, WL76);
sram_cell_6t_3 inst_cell_76_114 ( BL114, BLN114, WL76);
sram_cell_6t_3 inst_cell_76_113 ( BL113, BLN113, WL76);
sram_cell_6t_3 inst_cell_76_112 ( BL112, BLN112, WL76);
sram_cell_6t_3 inst_cell_76_111 ( BL111, BLN111, WL76);
sram_cell_6t_3 inst_cell_76_110 ( BL110, BLN110, WL76);
sram_cell_6t_3 inst_cell_76_109 ( BL109, BLN109, WL76);
sram_cell_6t_3 inst_cell_76_108 ( BL108, BLN108, WL76);
sram_cell_6t_3 inst_cell_76_107 ( BL107, BLN107, WL76);
sram_cell_6t_3 inst_cell_76_106 ( BL106, BLN106, WL76);
sram_cell_6t_3 inst_cell_76_105 ( BL105, BLN105, WL76);
sram_cell_6t_3 inst_cell_76_104 ( BL104, BLN104, WL76);
sram_cell_6t_3 inst_cell_76_103 ( BL103, BLN103, WL76);
sram_cell_6t_3 inst_cell_76_102 ( BL102, BLN102, WL76);
sram_cell_6t_3 inst_cell_76_101 ( BL101, BLN101, WL76);
sram_cell_6t_3 inst_cell_76_100 ( BL100, BLN100, WL76);
sram_cell_6t_3 inst_cell_76_99 ( BL99, BLN99, WL76);
sram_cell_6t_3 inst_cell_76_98 ( BL98, BLN98, WL76);
sram_cell_6t_3 inst_cell_76_97 ( BL97, BLN97, WL76);
sram_cell_6t_3 inst_cell_76_96 ( BL96, BLN96, WL76);
sram_cell_6t_3 inst_cell_76_95 ( BL95, BLN95, WL76);
sram_cell_6t_3 inst_cell_76_94 ( BL94, BLN94, WL76);
sram_cell_6t_3 inst_cell_76_93 ( BL93, BLN93, WL76);
sram_cell_6t_3 inst_cell_76_92 ( BL92, BLN92, WL76);
sram_cell_6t_3 inst_cell_76_91 ( BL91, BLN91, WL76);
sram_cell_6t_3 inst_cell_76_90 ( BL90, BLN90, WL76);
sram_cell_6t_3 inst_cell_76_89 ( BL89, BLN89, WL76);
sram_cell_6t_3 inst_cell_76_88 ( BL88, BLN88, WL76);
sram_cell_6t_3 inst_cell_76_87 ( BL87, BLN87, WL76);
sram_cell_6t_3 inst_cell_76_86 ( BL86, BLN86, WL76);
sram_cell_6t_3 inst_cell_76_85 ( BL85, BLN85, WL76);
sram_cell_6t_3 inst_cell_76_84 ( BL84, BLN84, WL76);
sram_cell_6t_3 inst_cell_76_83 ( BL83, BLN83, WL76);
sram_cell_6t_3 inst_cell_76_82 ( BL82, BLN82, WL76);
sram_cell_6t_3 inst_cell_76_81 ( BL81, BLN81, WL76);
sram_cell_6t_3 inst_cell_76_80 ( BL80, BLN80, WL76);
sram_cell_6t_3 inst_cell_76_79 ( BL79, BLN79, WL76);
sram_cell_6t_3 inst_cell_76_78 ( BL78, BLN78, WL76);
sram_cell_6t_3 inst_cell_76_77 ( BL77, BLN77, WL76);
sram_cell_6t_3 inst_cell_76_76 ( BL76, BLN76, WL76);
sram_cell_6t_3 inst_cell_76_75 ( BL75, BLN75, WL76);
sram_cell_6t_3 inst_cell_76_74 ( BL74, BLN74, WL76);
sram_cell_6t_3 inst_cell_76_73 ( BL73, BLN73, WL76);
sram_cell_6t_3 inst_cell_76_72 ( BL72, BLN72, WL76);
sram_cell_6t_3 inst_cell_76_71 ( BL71, BLN71, WL76);
sram_cell_6t_3 inst_cell_76_70 ( BL70, BLN70, WL76);
sram_cell_6t_3 inst_cell_76_69 ( BL69, BLN69, WL76);
sram_cell_6t_3 inst_cell_76_68 ( BL68, BLN68, WL76);
sram_cell_6t_3 inst_cell_76_67 ( BL67, BLN67, WL76);
sram_cell_6t_3 inst_cell_76_66 ( BL66, BLN66, WL76);
sram_cell_6t_3 inst_cell_76_65 ( BL65, BLN65, WL76);
sram_cell_6t_3 inst_cell_76_64 ( BL64, BLN64, WL76);
sram_cell_6t_3 inst_cell_76_63 ( BL63, BLN63, WL76);
sram_cell_6t_3 inst_cell_76_62 ( BL62, BLN62, WL76);
sram_cell_6t_3 inst_cell_76_61 ( BL61, BLN61, WL76);
sram_cell_6t_3 inst_cell_76_60 ( BL60, BLN60, WL76);
sram_cell_6t_3 inst_cell_76_59 ( BL59, BLN59, WL76);
sram_cell_6t_3 inst_cell_76_58 ( BL58, BLN58, WL76);
sram_cell_6t_3 inst_cell_76_57 ( BL57, BLN57, WL76);
sram_cell_6t_3 inst_cell_76_56 ( BL56, BLN56, WL76);
sram_cell_6t_3 inst_cell_76_55 ( BL55, BLN55, WL76);
sram_cell_6t_3 inst_cell_76_54 ( BL54, BLN54, WL76);
sram_cell_6t_3 inst_cell_76_53 ( BL53, BLN53, WL76);
sram_cell_6t_3 inst_cell_76_52 ( BL52, BLN52, WL76);
sram_cell_6t_3 inst_cell_76_51 ( BL51, BLN51, WL76);
sram_cell_6t_3 inst_cell_76_50 ( BL50, BLN50, WL76);
sram_cell_6t_3 inst_cell_76_49 ( BL49, BLN49, WL76);
sram_cell_6t_3 inst_cell_76_48 ( BL48, BLN48, WL76);
sram_cell_6t_3 inst_cell_76_47 ( BL47, BLN47, WL76);
sram_cell_6t_3 inst_cell_76_46 ( BL46, BLN46, WL76);
sram_cell_6t_3 inst_cell_76_45 ( BL45, BLN45, WL76);
sram_cell_6t_3 inst_cell_76_44 ( BL44, BLN44, WL76);
sram_cell_6t_3 inst_cell_76_43 ( BL43, BLN43, WL76);
sram_cell_6t_3 inst_cell_76_42 ( BL42, BLN42, WL76);
sram_cell_6t_3 inst_cell_76_41 ( BL41, BLN41, WL76);
sram_cell_6t_3 inst_cell_76_40 ( BL40, BLN40, WL76);
sram_cell_6t_3 inst_cell_76_39 ( BL39, BLN39, WL76);
sram_cell_6t_3 inst_cell_76_38 ( BL38, BLN38, WL76);
sram_cell_6t_3 inst_cell_76_37 ( BL37, BLN37, WL76);
sram_cell_6t_3 inst_cell_76_36 ( BL36, BLN36, WL76);
sram_cell_6t_3 inst_cell_76_35 ( BL35, BLN35, WL76);
sram_cell_6t_3 inst_cell_76_34 ( BL34, BLN34, WL76);
sram_cell_6t_3 inst_cell_76_33 ( BL33, BLN33, WL76);
sram_cell_6t_3 inst_cell_76_32 ( BL32, BLN32, WL76);
sram_cell_6t_3 inst_cell_76_31 ( BL31, BLN31, WL76);
sram_cell_6t_3 inst_cell_76_30 ( BL30, BLN30, WL76);
sram_cell_6t_3 inst_cell_76_29 ( BL29, BLN29, WL76);
sram_cell_6t_3 inst_cell_76_28 ( BL28, BLN28, WL76);
sram_cell_6t_3 inst_cell_76_27 ( BL27, BLN27, WL76);
sram_cell_6t_3 inst_cell_76_26 ( BL26, BLN26, WL76);
sram_cell_6t_3 inst_cell_76_25 ( BL25, BLN25, WL76);
sram_cell_6t_3 inst_cell_76_24 ( BL24, BLN24, WL76);
sram_cell_6t_3 inst_cell_76_23 ( BL23, BLN23, WL76);
sram_cell_6t_3 inst_cell_76_22 ( BL22, BLN22, WL76);
sram_cell_6t_3 inst_cell_76_21 ( BL21, BLN21, WL76);
sram_cell_6t_3 inst_cell_76_20 ( BL20, BLN20, WL76);
sram_cell_6t_3 inst_cell_76_19 ( BL19, BLN19, WL76);
sram_cell_6t_3 inst_cell_76_18 ( BL18, BLN18, WL76);
sram_cell_6t_3 inst_cell_76_17 ( BL17, BLN17, WL76);
sram_cell_6t_3 inst_cell_76_16 ( BL16, BLN16, WL76);
sram_cell_6t_3 inst_cell_76_15 ( BL15, BLN15, WL76);
sram_cell_6t_3 inst_cell_76_14 ( BL14, BLN14, WL76);
sram_cell_6t_3 inst_cell_76_13 ( BL13, BLN13, WL76);
sram_cell_6t_3 inst_cell_76_12 ( BL12, BLN12, WL76);
sram_cell_6t_3 inst_cell_76_11 ( BL11, BLN11, WL76);
sram_cell_6t_3 inst_cell_76_10 ( BL10, BLN10, WL76);
sram_cell_6t_3 inst_cell_76_9 ( BL9, BLN9, WL76);
sram_cell_6t_3 inst_cell_76_8 ( BL8, BLN8, WL76);
sram_cell_6t_3 inst_cell_76_7 ( BL7, BLN7, WL76);
sram_cell_6t_3 inst_cell_76_6 ( BL6, BLN6, WL76);
sram_cell_6t_3 inst_cell_76_5 ( BL5, BLN5, WL76);
sram_cell_6t_3 inst_cell_76_4 ( BL4, BLN4, WL76);
sram_cell_6t_3 inst_cell_76_3 ( BL3, BLN3, WL76);
sram_cell_6t_3 inst_cell_76_2 ( BL2, BLN2, WL76);
sram_cell_6t_3 inst_cell_76_1 ( BL1, BLN1, WL76);
sram_cell_6t_3 inst_cell_76_0 ( BL0, BLN0, WL76);
sram_cell_6t_3 inst_cell_75_127 ( BL127, BLN127, WL75);
sram_cell_6t_3 inst_cell_75_126 ( BL126, BLN126, WL75);
sram_cell_6t_3 inst_cell_75_125 ( BL125, BLN125, WL75);
sram_cell_6t_3 inst_cell_75_124 ( BL124, BLN124, WL75);
sram_cell_6t_3 inst_cell_75_123 ( BL123, BLN123, WL75);
sram_cell_6t_3 inst_cell_75_122 ( BL122, BLN122, WL75);
sram_cell_6t_3 inst_cell_75_121 ( BL121, BLN121, WL75);
sram_cell_6t_3 inst_cell_75_120 ( BL120, BLN120, WL75);
sram_cell_6t_3 inst_cell_75_119 ( BL119, BLN119, WL75);
sram_cell_6t_3 inst_cell_75_118 ( BL118, BLN118, WL75);
sram_cell_6t_3 inst_cell_75_117 ( BL117, BLN117, WL75);
sram_cell_6t_3 inst_cell_75_116 ( BL116, BLN116, WL75);
sram_cell_6t_3 inst_cell_75_115 ( BL115, BLN115, WL75);
sram_cell_6t_3 inst_cell_75_114 ( BL114, BLN114, WL75);
sram_cell_6t_3 inst_cell_75_113 ( BL113, BLN113, WL75);
sram_cell_6t_3 inst_cell_75_112 ( BL112, BLN112, WL75);
sram_cell_6t_3 inst_cell_75_111 ( BL111, BLN111, WL75);
sram_cell_6t_3 inst_cell_75_110 ( BL110, BLN110, WL75);
sram_cell_6t_3 inst_cell_75_109 ( BL109, BLN109, WL75);
sram_cell_6t_3 inst_cell_75_108 ( BL108, BLN108, WL75);
sram_cell_6t_3 inst_cell_75_107 ( BL107, BLN107, WL75);
sram_cell_6t_3 inst_cell_75_106 ( BL106, BLN106, WL75);
sram_cell_6t_3 inst_cell_75_105 ( BL105, BLN105, WL75);
sram_cell_6t_3 inst_cell_75_104 ( BL104, BLN104, WL75);
sram_cell_6t_3 inst_cell_75_103 ( BL103, BLN103, WL75);
sram_cell_6t_3 inst_cell_75_102 ( BL102, BLN102, WL75);
sram_cell_6t_3 inst_cell_75_101 ( BL101, BLN101, WL75);
sram_cell_6t_3 inst_cell_75_100 ( BL100, BLN100, WL75);
sram_cell_6t_3 inst_cell_75_99 ( BL99, BLN99, WL75);
sram_cell_6t_3 inst_cell_75_98 ( BL98, BLN98, WL75);
sram_cell_6t_3 inst_cell_75_97 ( BL97, BLN97, WL75);
sram_cell_6t_3 inst_cell_75_96 ( BL96, BLN96, WL75);
sram_cell_6t_3 inst_cell_75_95 ( BL95, BLN95, WL75);
sram_cell_6t_3 inst_cell_75_94 ( BL94, BLN94, WL75);
sram_cell_6t_3 inst_cell_75_93 ( BL93, BLN93, WL75);
sram_cell_6t_3 inst_cell_75_92 ( BL92, BLN92, WL75);
sram_cell_6t_3 inst_cell_75_91 ( BL91, BLN91, WL75);
sram_cell_6t_3 inst_cell_75_90 ( BL90, BLN90, WL75);
sram_cell_6t_3 inst_cell_75_89 ( BL89, BLN89, WL75);
sram_cell_6t_3 inst_cell_75_88 ( BL88, BLN88, WL75);
sram_cell_6t_3 inst_cell_75_87 ( BL87, BLN87, WL75);
sram_cell_6t_3 inst_cell_75_86 ( BL86, BLN86, WL75);
sram_cell_6t_3 inst_cell_75_85 ( BL85, BLN85, WL75);
sram_cell_6t_3 inst_cell_75_84 ( BL84, BLN84, WL75);
sram_cell_6t_3 inst_cell_75_83 ( BL83, BLN83, WL75);
sram_cell_6t_3 inst_cell_75_82 ( BL82, BLN82, WL75);
sram_cell_6t_3 inst_cell_75_81 ( BL81, BLN81, WL75);
sram_cell_6t_3 inst_cell_75_80 ( BL80, BLN80, WL75);
sram_cell_6t_3 inst_cell_75_79 ( BL79, BLN79, WL75);
sram_cell_6t_3 inst_cell_75_78 ( BL78, BLN78, WL75);
sram_cell_6t_3 inst_cell_75_77 ( BL77, BLN77, WL75);
sram_cell_6t_3 inst_cell_75_76 ( BL76, BLN76, WL75);
sram_cell_6t_3 inst_cell_75_75 ( BL75, BLN75, WL75);
sram_cell_6t_3 inst_cell_75_74 ( BL74, BLN74, WL75);
sram_cell_6t_3 inst_cell_75_73 ( BL73, BLN73, WL75);
sram_cell_6t_3 inst_cell_75_72 ( BL72, BLN72, WL75);
sram_cell_6t_3 inst_cell_75_71 ( BL71, BLN71, WL75);
sram_cell_6t_3 inst_cell_75_70 ( BL70, BLN70, WL75);
sram_cell_6t_3 inst_cell_75_69 ( BL69, BLN69, WL75);
sram_cell_6t_3 inst_cell_75_68 ( BL68, BLN68, WL75);
sram_cell_6t_3 inst_cell_75_67 ( BL67, BLN67, WL75);
sram_cell_6t_3 inst_cell_75_66 ( BL66, BLN66, WL75);
sram_cell_6t_3 inst_cell_75_65 ( BL65, BLN65, WL75);
sram_cell_6t_3 inst_cell_75_64 ( BL64, BLN64, WL75);
sram_cell_6t_3 inst_cell_75_63 ( BL63, BLN63, WL75);
sram_cell_6t_3 inst_cell_75_62 ( BL62, BLN62, WL75);
sram_cell_6t_3 inst_cell_75_61 ( BL61, BLN61, WL75);
sram_cell_6t_3 inst_cell_75_60 ( BL60, BLN60, WL75);
sram_cell_6t_3 inst_cell_75_59 ( BL59, BLN59, WL75);
sram_cell_6t_3 inst_cell_75_58 ( BL58, BLN58, WL75);
sram_cell_6t_3 inst_cell_75_57 ( BL57, BLN57, WL75);
sram_cell_6t_3 inst_cell_75_56 ( BL56, BLN56, WL75);
sram_cell_6t_3 inst_cell_75_55 ( BL55, BLN55, WL75);
sram_cell_6t_3 inst_cell_75_54 ( BL54, BLN54, WL75);
sram_cell_6t_3 inst_cell_75_53 ( BL53, BLN53, WL75);
sram_cell_6t_3 inst_cell_75_52 ( BL52, BLN52, WL75);
sram_cell_6t_3 inst_cell_75_51 ( BL51, BLN51, WL75);
sram_cell_6t_3 inst_cell_75_50 ( BL50, BLN50, WL75);
sram_cell_6t_3 inst_cell_75_49 ( BL49, BLN49, WL75);
sram_cell_6t_3 inst_cell_75_48 ( BL48, BLN48, WL75);
sram_cell_6t_3 inst_cell_75_47 ( BL47, BLN47, WL75);
sram_cell_6t_3 inst_cell_75_46 ( BL46, BLN46, WL75);
sram_cell_6t_3 inst_cell_75_45 ( BL45, BLN45, WL75);
sram_cell_6t_3 inst_cell_75_44 ( BL44, BLN44, WL75);
sram_cell_6t_3 inst_cell_75_43 ( BL43, BLN43, WL75);
sram_cell_6t_3 inst_cell_75_42 ( BL42, BLN42, WL75);
sram_cell_6t_3 inst_cell_75_41 ( BL41, BLN41, WL75);
sram_cell_6t_3 inst_cell_75_40 ( BL40, BLN40, WL75);
sram_cell_6t_3 inst_cell_75_39 ( BL39, BLN39, WL75);
sram_cell_6t_3 inst_cell_75_38 ( BL38, BLN38, WL75);
sram_cell_6t_3 inst_cell_75_37 ( BL37, BLN37, WL75);
sram_cell_6t_3 inst_cell_75_36 ( BL36, BLN36, WL75);
sram_cell_6t_3 inst_cell_75_35 ( BL35, BLN35, WL75);
sram_cell_6t_3 inst_cell_75_34 ( BL34, BLN34, WL75);
sram_cell_6t_3 inst_cell_75_33 ( BL33, BLN33, WL75);
sram_cell_6t_3 inst_cell_75_32 ( BL32, BLN32, WL75);
sram_cell_6t_3 inst_cell_75_31 ( BL31, BLN31, WL75);
sram_cell_6t_3 inst_cell_75_30 ( BL30, BLN30, WL75);
sram_cell_6t_3 inst_cell_75_29 ( BL29, BLN29, WL75);
sram_cell_6t_3 inst_cell_75_28 ( BL28, BLN28, WL75);
sram_cell_6t_3 inst_cell_75_27 ( BL27, BLN27, WL75);
sram_cell_6t_3 inst_cell_75_26 ( BL26, BLN26, WL75);
sram_cell_6t_3 inst_cell_75_25 ( BL25, BLN25, WL75);
sram_cell_6t_3 inst_cell_75_24 ( BL24, BLN24, WL75);
sram_cell_6t_3 inst_cell_75_23 ( BL23, BLN23, WL75);
sram_cell_6t_3 inst_cell_75_22 ( BL22, BLN22, WL75);
sram_cell_6t_3 inst_cell_75_21 ( BL21, BLN21, WL75);
sram_cell_6t_3 inst_cell_75_20 ( BL20, BLN20, WL75);
sram_cell_6t_3 inst_cell_75_19 ( BL19, BLN19, WL75);
sram_cell_6t_3 inst_cell_75_18 ( BL18, BLN18, WL75);
sram_cell_6t_3 inst_cell_75_17 ( BL17, BLN17, WL75);
sram_cell_6t_3 inst_cell_75_16 ( BL16, BLN16, WL75);
sram_cell_6t_3 inst_cell_75_15 ( BL15, BLN15, WL75);
sram_cell_6t_3 inst_cell_75_14 ( BL14, BLN14, WL75);
sram_cell_6t_3 inst_cell_75_13 ( BL13, BLN13, WL75);
sram_cell_6t_3 inst_cell_75_12 ( BL12, BLN12, WL75);
sram_cell_6t_3 inst_cell_75_11 ( BL11, BLN11, WL75);
sram_cell_6t_3 inst_cell_75_10 ( BL10, BLN10, WL75);
sram_cell_6t_3 inst_cell_75_9 ( BL9, BLN9, WL75);
sram_cell_6t_3 inst_cell_75_8 ( BL8, BLN8, WL75);
sram_cell_6t_3 inst_cell_75_7 ( BL7, BLN7, WL75);
sram_cell_6t_3 inst_cell_75_6 ( BL6, BLN6, WL75);
sram_cell_6t_3 inst_cell_75_5 ( BL5, BLN5, WL75);
sram_cell_6t_3 inst_cell_75_4 ( BL4, BLN4, WL75);
sram_cell_6t_3 inst_cell_75_3 ( BL3, BLN3, WL75);
sram_cell_6t_3 inst_cell_75_2 ( BL2, BLN2, WL75);
sram_cell_6t_3 inst_cell_75_1 ( BL1, BLN1, WL75);
sram_cell_6t_3 inst_cell_75_0 ( BL0, BLN0, WL75);
sram_cell_6t_3 inst_cell_74_127 ( BL127, BLN127, WL74);
sram_cell_6t_3 inst_cell_74_126 ( BL126, BLN126, WL74);
sram_cell_6t_3 inst_cell_74_125 ( BL125, BLN125, WL74);
sram_cell_6t_3 inst_cell_74_124 ( BL124, BLN124, WL74);
sram_cell_6t_3 inst_cell_74_123 ( BL123, BLN123, WL74);
sram_cell_6t_3 inst_cell_74_122 ( BL122, BLN122, WL74);
sram_cell_6t_3 inst_cell_74_121 ( BL121, BLN121, WL74);
sram_cell_6t_3 inst_cell_74_120 ( BL120, BLN120, WL74);
sram_cell_6t_3 inst_cell_74_119 ( BL119, BLN119, WL74);
sram_cell_6t_3 inst_cell_74_118 ( BL118, BLN118, WL74);
sram_cell_6t_3 inst_cell_74_117 ( BL117, BLN117, WL74);
sram_cell_6t_3 inst_cell_74_116 ( BL116, BLN116, WL74);
sram_cell_6t_3 inst_cell_74_115 ( BL115, BLN115, WL74);
sram_cell_6t_3 inst_cell_74_114 ( BL114, BLN114, WL74);
sram_cell_6t_3 inst_cell_74_113 ( BL113, BLN113, WL74);
sram_cell_6t_3 inst_cell_74_112 ( BL112, BLN112, WL74);
sram_cell_6t_3 inst_cell_74_111 ( BL111, BLN111, WL74);
sram_cell_6t_3 inst_cell_74_110 ( BL110, BLN110, WL74);
sram_cell_6t_3 inst_cell_74_109 ( BL109, BLN109, WL74);
sram_cell_6t_3 inst_cell_74_108 ( BL108, BLN108, WL74);
sram_cell_6t_3 inst_cell_74_107 ( BL107, BLN107, WL74);
sram_cell_6t_3 inst_cell_74_106 ( BL106, BLN106, WL74);
sram_cell_6t_3 inst_cell_74_105 ( BL105, BLN105, WL74);
sram_cell_6t_3 inst_cell_74_104 ( BL104, BLN104, WL74);
sram_cell_6t_3 inst_cell_74_103 ( BL103, BLN103, WL74);
sram_cell_6t_3 inst_cell_74_102 ( BL102, BLN102, WL74);
sram_cell_6t_3 inst_cell_74_101 ( BL101, BLN101, WL74);
sram_cell_6t_3 inst_cell_74_100 ( BL100, BLN100, WL74);
sram_cell_6t_3 inst_cell_74_99 ( BL99, BLN99, WL74);
sram_cell_6t_3 inst_cell_74_98 ( BL98, BLN98, WL74);
sram_cell_6t_3 inst_cell_74_97 ( BL97, BLN97, WL74);
sram_cell_6t_3 inst_cell_74_96 ( BL96, BLN96, WL74);
sram_cell_6t_3 inst_cell_74_95 ( BL95, BLN95, WL74);
sram_cell_6t_3 inst_cell_74_94 ( BL94, BLN94, WL74);
sram_cell_6t_3 inst_cell_74_93 ( BL93, BLN93, WL74);
sram_cell_6t_3 inst_cell_74_92 ( BL92, BLN92, WL74);
sram_cell_6t_3 inst_cell_74_91 ( BL91, BLN91, WL74);
sram_cell_6t_3 inst_cell_74_90 ( BL90, BLN90, WL74);
sram_cell_6t_3 inst_cell_74_89 ( BL89, BLN89, WL74);
sram_cell_6t_3 inst_cell_74_88 ( BL88, BLN88, WL74);
sram_cell_6t_3 inst_cell_74_87 ( BL87, BLN87, WL74);
sram_cell_6t_3 inst_cell_74_86 ( BL86, BLN86, WL74);
sram_cell_6t_3 inst_cell_74_85 ( BL85, BLN85, WL74);
sram_cell_6t_3 inst_cell_74_84 ( BL84, BLN84, WL74);
sram_cell_6t_3 inst_cell_74_83 ( BL83, BLN83, WL74);
sram_cell_6t_3 inst_cell_74_82 ( BL82, BLN82, WL74);
sram_cell_6t_3 inst_cell_74_81 ( BL81, BLN81, WL74);
sram_cell_6t_3 inst_cell_74_80 ( BL80, BLN80, WL74);
sram_cell_6t_3 inst_cell_74_79 ( BL79, BLN79, WL74);
sram_cell_6t_3 inst_cell_74_78 ( BL78, BLN78, WL74);
sram_cell_6t_3 inst_cell_74_77 ( BL77, BLN77, WL74);
sram_cell_6t_3 inst_cell_74_76 ( BL76, BLN76, WL74);
sram_cell_6t_3 inst_cell_74_75 ( BL75, BLN75, WL74);
sram_cell_6t_3 inst_cell_74_74 ( BL74, BLN74, WL74);
sram_cell_6t_3 inst_cell_74_73 ( BL73, BLN73, WL74);
sram_cell_6t_3 inst_cell_74_72 ( BL72, BLN72, WL74);
sram_cell_6t_3 inst_cell_74_71 ( BL71, BLN71, WL74);
sram_cell_6t_3 inst_cell_74_70 ( BL70, BLN70, WL74);
sram_cell_6t_3 inst_cell_74_69 ( BL69, BLN69, WL74);
sram_cell_6t_3 inst_cell_74_68 ( BL68, BLN68, WL74);
sram_cell_6t_3 inst_cell_74_67 ( BL67, BLN67, WL74);
sram_cell_6t_3 inst_cell_74_66 ( BL66, BLN66, WL74);
sram_cell_6t_3 inst_cell_74_65 ( BL65, BLN65, WL74);
sram_cell_6t_3 inst_cell_74_64 ( BL64, BLN64, WL74);
sram_cell_6t_3 inst_cell_74_63 ( BL63, BLN63, WL74);
sram_cell_6t_3 inst_cell_74_62 ( BL62, BLN62, WL74);
sram_cell_6t_3 inst_cell_74_61 ( BL61, BLN61, WL74);
sram_cell_6t_3 inst_cell_74_60 ( BL60, BLN60, WL74);
sram_cell_6t_3 inst_cell_74_59 ( BL59, BLN59, WL74);
sram_cell_6t_3 inst_cell_74_58 ( BL58, BLN58, WL74);
sram_cell_6t_3 inst_cell_74_57 ( BL57, BLN57, WL74);
sram_cell_6t_3 inst_cell_74_56 ( BL56, BLN56, WL74);
sram_cell_6t_3 inst_cell_74_55 ( BL55, BLN55, WL74);
sram_cell_6t_3 inst_cell_74_54 ( BL54, BLN54, WL74);
sram_cell_6t_3 inst_cell_74_53 ( BL53, BLN53, WL74);
sram_cell_6t_3 inst_cell_74_52 ( BL52, BLN52, WL74);
sram_cell_6t_3 inst_cell_74_51 ( BL51, BLN51, WL74);
sram_cell_6t_3 inst_cell_74_50 ( BL50, BLN50, WL74);
sram_cell_6t_3 inst_cell_74_49 ( BL49, BLN49, WL74);
sram_cell_6t_3 inst_cell_74_48 ( BL48, BLN48, WL74);
sram_cell_6t_3 inst_cell_74_47 ( BL47, BLN47, WL74);
sram_cell_6t_3 inst_cell_74_46 ( BL46, BLN46, WL74);
sram_cell_6t_3 inst_cell_74_45 ( BL45, BLN45, WL74);
sram_cell_6t_3 inst_cell_74_44 ( BL44, BLN44, WL74);
sram_cell_6t_3 inst_cell_74_43 ( BL43, BLN43, WL74);
sram_cell_6t_3 inst_cell_74_42 ( BL42, BLN42, WL74);
sram_cell_6t_3 inst_cell_74_41 ( BL41, BLN41, WL74);
sram_cell_6t_3 inst_cell_74_40 ( BL40, BLN40, WL74);
sram_cell_6t_3 inst_cell_74_39 ( BL39, BLN39, WL74);
sram_cell_6t_3 inst_cell_74_38 ( BL38, BLN38, WL74);
sram_cell_6t_3 inst_cell_74_37 ( BL37, BLN37, WL74);
sram_cell_6t_3 inst_cell_74_36 ( BL36, BLN36, WL74);
sram_cell_6t_3 inst_cell_74_35 ( BL35, BLN35, WL74);
sram_cell_6t_3 inst_cell_74_34 ( BL34, BLN34, WL74);
sram_cell_6t_3 inst_cell_74_33 ( BL33, BLN33, WL74);
sram_cell_6t_3 inst_cell_74_32 ( BL32, BLN32, WL74);
sram_cell_6t_3 inst_cell_74_31 ( BL31, BLN31, WL74);
sram_cell_6t_3 inst_cell_74_30 ( BL30, BLN30, WL74);
sram_cell_6t_3 inst_cell_74_29 ( BL29, BLN29, WL74);
sram_cell_6t_3 inst_cell_74_28 ( BL28, BLN28, WL74);
sram_cell_6t_3 inst_cell_74_27 ( BL27, BLN27, WL74);
sram_cell_6t_3 inst_cell_74_26 ( BL26, BLN26, WL74);
sram_cell_6t_3 inst_cell_74_25 ( BL25, BLN25, WL74);
sram_cell_6t_3 inst_cell_74_24 ( BL24, BLN24, WL74);
sram_cell_6t_3 inst_cell_74_23 ( BL23, BLN23, WL74);
sram_cell_6t_3 inst_cell_74_22 ( BL22, BLN22, WL74);
sram_cell_6t_3 inst_cell_74_21 ( BL21, BLN21, WL74);
sram_cell_6t_3 inst_cell_74_20 ( BL20, BLN20, WL74);
sram_cell_6t_3 inst_cell_74_19 ( BL19, BLN19, WL74);
sram_cell_6t_3 inst_cell_74_18 ( BL18, BLN18, WL74);
sram_cell_6t_3 inst_cell_74_17 ( BL17, BLN17, WL74);
sram_cell_6t_3 inst_cell_74_16 ( BL16, BLN16, WL74);
sram_cell_6t_3 inst_cell_74_15 ( BL15, BLN15, WL74);
sram_cell_6t_3 inst_cell_74_14 ( BL14, BLN14, WL74);
sram_cell_6t_3 inst_cell_74_13 ( BL13, BLN13, WL74);
sram_cell_6t_3 inst_cell_74_12 ( BL12, BLN12, WL74);
sram_cell_6t_3 inst_cell_74_11 ( BL11, BLN11, WL74);
sram_cell_6t_3 inst_cell_74_10 ( BL10, BLN10, WL74);
sram_cell_6t_3 inst_cell_74_9 ( BL9, BLN9, WL74);
sram_cell_6t_3 inst_cell_74_8 ( BL8, BLN8, WL74);
sram_cell_6t_3 inst_cell_74_7 ( BL7, BLN7, WL74);
sram_cell_6t_3 inst_cell_74_6 ( BL6, BLN6, WL74);
sram_cell_6t_3 inst_cell_74_5 ( BL5, BLN5, WL74);
sram_cell_6t_3 inst_cell_74_4 ( BL4, BLN4, WL74);
sram_cell_6t_3 inst_cell_74_3 ( BL3, BLN3, WL74);
sram_cell_6t_3 inst_cell_74_2 ( BL2, BLN2, WL74);
sram_cell_6t_3 inst_cell_74_1 ( BL1, BLN1, WL74);
sram_cell_6t_3 inst_cell_74_0 ( BL0, BLN0, WL74);
sram_cell_6t_3 inst_cell_73_127 ( BL127, BLN127, WL73);
sram_cell_6t_3 inst_cell_73_126 ( BL126, BLN126, WL73);
sram_cell_6t_3 inst_cell_73_125 ( BL125, BLN125, WL73);
sram_cell_6t_3 inst_cell_73_124 ( BL124, BLN124, WL73);
sram_cell_6t_3 inst_cell_73_123 ( BL123, BLN123, WL73);
sram_cell_6t_3 inst_cell_73_122 ( BL122, BLN122, WL73);
sram_cell_6t_3 inst_cell_73_121 ( BL121, BLN121, WL73);
sram_cell_6t_3 inst_cell_73_120 ( BL120, BLN120, WL73);
sram_cell_6t_3 inst_cell_73_119 ( BL119, BLN119, WL73);
sram_cell_6t_3 inst_cell_73_118 ( BL118, BLN118, WL73);
sram_cell_6t_3 inst_cell_73_117 ( BL117, BLN117, WL73);
sram_cell_6t_3 inst_cell_73_116 ( BL116, BLN116, WL73);
sram_cell_6t_3 inst_cell_73_115 ( BL115, BLN115, WL73);
sram_cell_6t_3 inst_cell_73_114 ( BL114, BLN114, WL73);
sram_cell_6t_3 inst_cell_73_113 ( BL113, BLN113, WL73);
sram_cell_6t_3 inst_cell_73_112 ( BL112, BLN112, WL73);
sram_cell_6t_3 inst_cell_73_111 ( BL111, BLN111, WL73);
sram_cell_6t_3 inst_cell_73_110 ( BL110, BLN110, WL73);
sram_cell_6t_3 inst_cell_73_109 ( BL109, BLN109, WL73);
sram_cell_6t_3 inst_cell_73_108 ( BL108, BLN108, WL73);
sram_cell_6t_3 inst_cell_73_107 ( BL107, BLN107, WL73);
sram_cell_6t_3 inst_cell_73_106 ( BL106, BLN106, WL73);
sram_cell_6t_3 inst_cell_73_105 ( BL105, BLN105, WL73);
sram_cell_6t_3 inst_cell_73_104 ( BL104, BLN104, WL73);
sram_cell_6t_3 inst_cell_73_103 ( BL103, BLN103, WL73);
sram_cell_6t_3 inst_cell_73_102 ( BL102, BLN102, WL73);
sram_cell_6t_3 inst_cell_73_101 ( BL101, BLN101, WL73);
sram_cell_6t_3 inst_cell_73_100 ( BL100, BLN100, WL73);
sram_cell_6t_3 inst_cell_73_99 ( BL99, BLN99, WL73);
sram_cell_6t_3 inst_cell_73_98 ( BL98, BLN98, WL73);
sram_cell_6t_3 inst_cell_73_97 ( BL97, BLN97, WL73);
sram_cell_6t_3 inst_cell_73_96 ( BL96, BLN96, WL73);
sram_cell_6t_3 inst_cell_73_95 ( BL95, BLN95, WL73);
sram_cell_6t_3 inst_cell_73_94 ( BL94, BLN94, WL73);
sram_cell_6t_3 inst_cell_73_93 ( BL93, BLN93, WL73);
sram_cell_6t_3 inst_cell_73_92 ( BL92, BLN92, WL73);
sram_cell_6t_3 inst_cell_73_91 ( BL91, BLN91, WL73);
sram_cell_6t_3 inst_cell_73_90 ( BL90, BLN90, WL73);
sram_cell_6t_3 inst_cell_73_89 ( BL89, BLN89, WL73);
sram_cell_6t_3 inst_cell_73_88 ( BL88, BLN88, WL73);
sram_cell_6t_3 inst_cell_73_87 ( BL87, BLN87, WL73);
sram_cell_6t_3 inst_cell_73_86 ( BL86, BLN86, WL73);
sram_cell_6t_3 inst_cell_73_85 ( BL85, BLN85, WL73);
sram_cell_6t_3 inst_cell_73_84 ( BL84, BLN84, WL73);
sram_cell_6t_3 inst_cell_73_83 ( BL83, BLN83, WL73);
sram_cell_6t_3 inst_cell_73_82 ( BL82, BLN82, WL73);
sram_cell_6t_3 inst_cell_73_81 ( BL81, BLN81, WL73);
sram_cell_6t_3 inst_cell_73_80 ( BL80, BLN80, WL73);
sram_cell_6t_3 inst_cell_73_79 ( BL79, BLN79, WL73);
sram_cell_6t_3 inst_cell_73_78 ( BL78, BLN78, WL73);
sram_cell_6t_3 inst_cell_73_77 ( BL77, BLN77, WL73);
sram_cell_6t_3 inst_cell_73_76 ( BL76, BLN76, WL73);
sram_cell_6t_3 inst_cell_73_75 ( BL75, BLN75, WL73);
sram_cell_6t_3 inst_cell_73_74 ( BL74, BLN74, WL73);
sram_cell_6t_3 inst_cell_73_73 ( BL73, BLN73, WL73);
sram_cell_6t_3 inst_cell_73_72 ( BL72, BLN72, WL73);
sram_cell_6t_3 inst_cell_73_71 ( BL71, BLN71, WL73);
sram_cell_6t_3 inst_cell_73_70 ( BL70, BLN70, WL73);
sram_cell_6t_3 inst_cell_73_69 ( BL69, BLN69, WL73);
sram_cell_6t_3 inst_cell_73_68 ( BL68, BLN68, WL73);
sram_cell_6t_3 inst_cell_73_67 ( BL67, BLN67, WL73);
sram_cell_6t_3 inst_cell_73_66 ( BL66, BLN66, WL73);
sram_cell_6t_3 inst_cell_73_65 ( BL65, BLN65, WL73);
sram_cell_6t_3 inst_cell_73_64 ( BL64, BLN64, WL73);
sram_cell_6t_3 inst_cell_73_63 ( BL63, BLN63, WL73);
sram_cell_6t_3 inst_cell_73_62 ( BL62, BLN62, WL73);
sram_cell_6t_3 inst_cell_73_61 ( BL61, BLN61, WL73);
sram_cell_6t_3 inst_cell_73_60 ( BL60, BLN60, WL73);
sram_cell_6t_3 inst_cell_73_59 ( BL59, BLN59, WL73);
sram_cell_6t_3 inst_cell_73_58 ( BL58, BLN58, WL73);
sram_cell_6t_3 inst_cell_73_57 ( BL57, BLN57, WL73);
sram_cell_6t_3 inst_cell_73_56 ( BL56, BLN56, WL73);
sram_cell_6t_3 inst_cell_73_55 ( BL55, BLN55, WL73);
sram_cell_6t_3 inst_cell_73_54 ( BL54, BLN54, WL73);
sram_cell_6t_3 inst_cell_73_53 ( BL53, BLN53, WL73);
sram_cell_6t_3 inst_cell_73_52 ( BL52, BLN52, WL73);
sram_cell_6t_3 inst_cell_73_51 ( BL51, BLN51, WL73);
sram_cell_6t_3 inst_cell_73_50 ( BL50, BLN50, WL73);
sram_cell_6t_3 inst_cell_73_49 ( BL49, BLN49, WL73);
sram_cell_6t_3 inst_cell_73_48 ( BL48, BLN48, WL73);
sram_cell_6t_3 inst_cell_73_47 ( BL47, BLN47, WL73);
sram_cell_6t_3 inst_cell_73_46 ( BL46, BLN46, WL73);
sram_cell_6t_3 inst_cell_73_45 ( BL45, BLN45, WL73);
sram_cell_6t_3 inst_cell_73_44 ( BL44, BLN44, WL73);
sram_cell_6t_3 inst_cell_73_43 ( BL43, BLN43, WL73);
sram_cell_6t_3 inst_cell_73_42 ( BL42, BLN42, WL73);
sram_cell_6t_3 inst_cell_73_41 ( BL41, BLN41, WL73);
sram_cell_6t_3 inst_cell_73_40 ( BL40, BLN40, WL73);
sram_cell_6t_3 inst_cell_73_39 ( BL39, BLN39, WL73);
sram_cell_6t_3 inst_cell_73_38 ( BL38, BLN38, WL73);
sram_cell_6t_3 inst_cell_73_37 ( BL37, BLN37, WL73);
sram_cell_6t_3 inst_cell_73_36 ( BL36, BLN36, WL73);
sram_cell_6t_3 inst_cell_73_35 ( BL35, BLN35, WL73);
sram_cell_6t_3 inst_cell_73_34 ( BL34, BLN34, WL73);
sram_cell_6t_3 inst_cell_73_33 ( BL33, BLN33, WL73);
sram_cell_6t_3 inst_cell_73_32 ( BL32, BLN32, WL73);
sram_cell_6t_3 inst_cell_73_31 ( BL31, BLN31, WL73);
sram_cell_6t_3 inst_cell_73_30 ( BL30, BLN30, WL73);
sram_cell_6t_3 inst_cell_73_29 ( BL29, BLN29, WL73);
sram_cell_6t_3 inst_cell_73_28 ( BL28, BLN28, WL73);
sram_cell_6t_3 inst_cell_73_27 ( BL27, BLN27, WL73);
sram_cell_6t_3 inst_cell_73_26 ( BL26, BLN26, WL73);
sram_cell_6t_3 inst_cell_73_25 ( BL25, BLN25, WL73);
sram_cell_6t_3 inst_cell_73_24 ( BL24, BLN24, WL73);
sram_cell_6t_3 inst_cell_73_23 ( BL23, BLN23, WL73);
sram_cell_6t_3 inst_cell_73_22 ( BL22, BLN22, WL73);
sram_cell_6t_3 inst_cell_73_21 ( BL21, BLN21, WL73);
sram_cell_6t_3 inst_cell_73_20 ( BL20, BLN20, WL73);
sram_cell_6t_3 inst_cell_73_19 ( BL19, BLN19, WL73);
sram_cell_6t_3 inst_cell_73_18 ( BL18, BLN18, WL73);
sram_cell_6t_3 inst_cell_73_17 ( BL17, BLN17, WL73);
sram_cell_6t_3 inst_cell_73_16 ( BL16, BLN16, WL73);
sram_cell_6t_3 inst_cell_73_15 ( BL15, BLN15, WL73);
sram_cell_6t_3 inst_cell_73_14 ( BL14, BLN14, WL73);
sram_cell_6t_3 inst_cell_73_13 ( BL13, BLN13, WL73);
sram_cell_6t_3 inst_cell_73_12 ( BL12, BLN12, WL73);
sram_cell_6t_3 inst_cell_73_11 ( BL11, BLN11, WL73);
sram_cell_6t_3 inst_cell_73_10 ( BL10, BLN10, WL73);
sram_cell_6t_3 inst_cell_73_9 ( BL9, BLN9, WL73);
sram_cell_6t_3 inst_cell_73_8 ( BL8, BLN8, WL73);
sram_cell_6t_3 inst_cell_73_7 ( BL7, BLN7, WL73);
sram_cell_6t_3 inst_cell_73_6 ( BL6, BLN6, WL73);
sram_cell_6t_3 inst_cell_73_5 ( BL5, BLN5, WL73);
sram_cell_6t_3 inst_cell_73_4 ( BL4, BLN4, WL73);
sram_cell_6t_3 inst_cell_73_3 ( BL3, BLN3, WL73);
sram_cell_6t_3 inst_cell_73_2 ( BL2, BLN2, WL73);
sram_cell_6t_3 inst_cell_73_1 ( BL1, BLN1, WL73);
sram_cell_6t_3 inst_cell_73_0 ( BL0, BLN0, WL73);
sram_cell_6t_3 inst_cell_72_127 ( BL127, BLN127, WL72);
sram_cell_6t_3 inst_cell_72_126 ( BL126, BLN126, WL72);
sram_cell_6t_3 inst_cell_72_125 ( BL125, BLN125, WL72);
sram_cell_6t_3 inst_cell_72_124 ( BL124, BLN124, WL72);
sram_cell_6t_3 inst_cell_72_123 ( BL123, BLN123, WL72);
sram_cell_6t_3 inst_cell_72_122 ( BL122, BLN122, WL72);
sram_cell_6t_3 inst_cell_72_121 ( BL121, BLN121, WL72);
sram_cell_6t_3 inst_cell_72_120 ( BL120, BLN120, WL72);
sram_cell_6t_3 inst_cell_72_119 ( BL119, BLN119, WL72);
sram_cell_6t_3 inst_cell_72_118 ( BL118, BLN118, WL72);
sram_cell_6t_3 inst_cell_72_117 ( BL117, BLN117, WL72);
sram_cell_6t_3 inst_cell_72_116 ( BL116, BLN116, WL72);
sram_cell_6t_3 inst_cell_72_115 ( BL115, BLN115, WL72);
sram_cell_6t_3 inst_cell_72_114 ( BL114, BLN114, WL72);
sram_cell_6t_3 inst_cell_72_113 ( BL113, BLN113, WL72);
sram_cell_6t_3 inst_cell_72_112 ( BL112, BLN112, WL72);
sram_cell_6t_3 inst_cell_72_111 ( BL111, BLN111, WL72);
sram_cell_6t_3 inst_cell_72_110 ( BL110, BLN110, WL72);
sram_cell_6t_3 inst_cell_72_109 ( BL109, BLN109, WL72);
sram_cell_6t_3 inst_cell_72_108 ( BL108, BLN108, WL72);
sram_cell_6t_3 inst_cell_72_107 ( BL107, BLN107, WL72);
sram_cell_6t_3 inst_cell_72_106 ( BL106, BLN106, WL72);
sram_cell_6t_3 inst_cell_72_105 ( BL105, BLN105, WL72);
sram_cell_6t_3 inst_cell_72_104 ( BL104, BLN104, WL72);
sram_cell_6t_3 inst_cell_72_103 ( BL103, BLN103, WL72);
sram_cell_6t_3 inst_cell_72_102 ( BL102, BLN102, WL72);
sram_cell_6t_3 inst_cell_72_101 ( BL101, BLN101, WL72);
sram_cell_6t_3 inst_cell_72_100 ( BL100, BLN100, WL72);
sram_cell_6t_3 inst_cell_72_99 ( BL99, BLN99, WL72);
sram_cell_6t_3 inst_cell_72_98 ( BL98, BLN98, WL72);
sram_cell_6t_3 inst_cell_72_97 ( BL97, BLN97, WL72);
sram_cell_6t_3 inst_cell_72_96 ( BL96, BLN96, WL72);
sram_cell_6t_3 inst_cell_72_95 ( BL95, BLN95, WL72);
sram_cell_6t_3 inst_cell_72_94 ( BL94, BLN94, WL72);
sram_cell_6t_3 inst_cell_72_93 ( BL93, BLN93, WL72);
sram_cell_6t_3 inst_cell_72_92 ( BL92, BLN92, WL72);
sram_cell_6t_3 inst_cell_72_91 ( BL91, BLN91, WL72);
sram_cell_6t_3 inst_cell_72_90 ( BL90, BLN90, WL72);
sram_cell_6t_3 inst_cell_72_89 ( BL89, BLN89, WL72);
sram_cell_6t_3 inst_cell_72_88 ( BL88, BLN88, WL72);
sram_cell_6t_3 inst_cell_72_87 ( BL87, BLN87, WL72);
sram_cell_6t_3 inst_cell_72_86 ( BL86, BLN86, WL72);
sram_cell_6t_3 inst_cell_72_85 ( BL85, BLN85, WL72);
sram_cell_6t_3 inst_cell_72_84 ( BL84, BLN84, WL72);
sram_cell_6t_3 inst_cell_72_83 ( BL83, BLN83, WL72);
sram_cell_6t_3 inst_cell_72_82 ( BL82, BLN82, WL72);
sram_cell_6t_3 inst_cell_72_81 ( BL81, BLN81, WL72);
sram_cell_6t_3 inst_cell_72_80 ( BL80, BLN80, WL72);
sram_cell_6t_3 inst_cell_72_79 ( BL79, BLN79, WL72);
sram_cell_6t_3 inst_cell_72_78 ( BL78, BLN78, WL72);
sram_cell_6t_3 inst_cell_72_77 ( BL77, BLN77, WL72);
sram_cell_6t_3 inst_cell_72_76 ( BL76, BLN76, WL72);
sram_cell_6t_3 inst_cell_72_75 ( BL75, BLN75, WL72);
sram_cell_6t_3 inst_cell_72_74 ( BL74, BLN74, WL72);
sram_cell_6t_3 inst_cell_72_73 ( BL73, BLN73, WL72);
sram_cell_6t_3 inst_cell_72_72 ( BL72, BLN72, WL72);
sram_cell_6t_3 inst_cell_72_71 ( BL71, BLN71, WL72);
sram_cell_6t_3 inst_cell_72_70 ( BL70, BLN70, WL72);
sram_cell_6t_3 inst_cell_72_69 ( BL69, BLN69, WL72);
sram_cell_6t_3 inst_cell_72_68 ( BL68, BLN68, WL72);
sram_cell_6t_3 inst_cell_72_67 ( BL67, BLN67, WL72);
sram_cell_6t_3 inst_cell_72_66 ( BL66, BLN66, WL72);
sram_cell_6t_3 inst_cell_72_65 ( BL65, BLN65, WL72);
sram_cell_6t_3 inst_cell_72_64 ( BL64, BLN64, WL72);
sram_cell_6t_3 inst_cell_72_63 ( BL63, BLN63, WL72);
sram_cell_6t_3 inst_cell_72_62 ( BL62, BLN62, WL72);
sram_cell_6t_3 inst_cell_72_61 ( BL61, BLN61, WL72);
sram_cell_6t_3 inst_cell_72_60 ( BL60, BLN60, WL72);
sram_cell_6t_3 inst_cell_72_59 ( BL59, BLN59, WL72);
sram_cell_6t_3 inst_cell_72_58 ( BL58, BLN58, WL72);
sram_cell_6t_3 inst_cell_72_57 ( BL57, BLN57, WL72);
sram_cell_6t_3 inst_cell_72_56 ( BL56, BLN56, WL72);
sram_cell_6t_3 inst_cell_72_55 ( BL55, BLN55, WL72);
sram_cell_6t_3 inst_cell_72_54 ( BL54, BLN54, WL72);
sram_cell_6t_3 inst_cell_72_53 ( BL53, BLN53, WL72);
sram_cell_6t_3 inst_cell_72_52 ( BL52, BLN52, WL72);
sram_cell_6t_3 inst_cell_72_51 ( BL51, BLN51, WL72);
sram_cell_6t_3 inst_cell_72_50 ( BL50, BLN50, WL72);
sram_cell_6t_3 inst_cell_72_49 ( BL49, BLN49, WL72);
sram_cell_6t_3 inst_cell_72_48 ( BL48, BLN48, WL72);
sram_cell_6t_3 inst_cell_72_47 ( BL47, BLN47, WL72);
sram_cell_6t_3 inst_cell_72_46 ( BL46, BLN46, WL72);
sram_cell_6t_3 inst_cell_72_45 ( BL45, BLN45, WL72);
sram_cell_6t_3 inst_cell_72_44 ( BL44, BLN44, WL72);
sram_cell_6t_3 inst_cell_72_43 ( BL43, BLN43, WL72);
sram_cell_6t_3 inst_cell_72_42 ( BL42, BLN42, WL72);
sram_cell_6t_3 inst_cell_72_41 ( BL41, BLN41, WL72);
sram_cell_6t_3 inst_cell_72_40 ( BL40, BLN40, WL72);
sram_cell_6t_3 inst_cell_72_39 ( BL39, BLN39, WL72);
sram_cell_6t_3 inst_cell_72_38 ( BL38, BLN38, WL72);
sram_cell_6t_3 inst_cell_72_37 ( BL37, BLN37, WL72);
sram_cell_6t_3 inst_cell_72_36 ( BL36, BLN36, WL72);
sram_cell_6t_3 inst_cell_72_35 ( BL35, BLN35, WL72);
sram_cell_6t_3 inst_cell_72_34 ( BL34, BLN34, WL72);
sram_cell_6t_3 inst_cell_72_33 ( BL33, BLN33, WL72);
sram_cell_6t_3 inst_cell_72_32 ( BL32, BLN32, WL72);
sram_cell_6t_3 inst_cell_72_31 ( BL31, BLN31, WL72);
sram_cell_6t_3 inst_cell_72_30 ( BL30, BLN30, WL72);
sram_cell_6t_3 inst_cell_72_29 ( BL29, BLN29, WL72);
sram_cell_6t_3 inst_cell_72_28 ( BL28, BLN28, WL72);
sram_cell_6t_3 inst_cell_72_27 ( BL27, BLN27, WL72);
sram_cell_6t_3 inst_cell_72_26 ( BL26, BLN26, WL72);
sram_cell_6t_3 inst_cell_72_25 ( BL25, BLN25, WL72);
sram_cell_6t_3 inst_cell_72_24 ( BL24, BLN24, WL72);
sram_cell_6t_3 inst_cell_72_23 ( BL23, BLN23, WL72);
sram_cell_6t_3 inst_cell_72_22 ( BL22, BLN22, WL72);
sram_cell_6t_3 inst_cell_72_21 ( BL21, BLN21, WL72);
sram_cell_6t_3 inst_cell_72_20 ( BL20, BLN20, WL72);
sram_cell_6t_3 inst_cell_72_19 ( BL19, BLN19, WL72);
sram_cell_6t_3 inst_cell_72_18 ( BL18, BLN18, WL72);
sram_cell_6t_3 inst_cell_72_17 ( BL17, BLN17, WL72);
sram_cell_6t_3 inst_cell_72_16 ( BL16, BLN16, WL72);
sram_cell_6t_3 inst_cell_72_15 ( BL15, BLN15, WL72);
sram_cell_6t_3 inst_cell_72_14 ( BL14, BLN14, WL72);
sram_cell_6t_3 inst_cell_72_13 ( BL13, BLN13, WL72);
sram_cell_6t_3 inst_cell_72_12 ( BL12, BLN12, WL72);
sram_cell_6t_3 inst_cell_72_11 ( BL11, BLN11, WL72);
sram_cell_6t_3 inst_cell_72_10 ( BL10, BLN10, WL72);
sram_cell_6t_3 inst_cell_72_9 ( BL9, BLN9, WL72);
sram_cell_6t_3 inst_cell_72_8 ( BL8, BLN8, WL72);
sram_cell_6t_3 inst_cell_72_7 ( BL7, BLN7, WL72);
sram_cell_6t_3 inst_cell_72_6 ( BL6, BLN6, WL72);
sram_cell_6t_3 inst_cell_72_5 ( BL5, BLN5, WL72);
sram_cell_6t_3 inst_cell_72_4 ( BL4, BLN4, WL72);
sram_cell_6t_3 inst_cell_72_3 ( BL3, BLN3, WL72);
sram_cell_6t_3 inst_cell_72_2 ( BL2, BLN2, WL72);
sram_cell_6t_3 inst_cell_72_1 ( BL1, BLN1, WL72);
sram_cell_6t_3 inst_cell_72_0 ( BL0, BLN0, WL72);
sram_cell_6t_3 inst_cell_71_127 ( BL127, BLN127, WL71);
sram_cell_6t_3 inst_cell_71_126 ( BL126, BLN126, WL71);
sram_cell_6t_3 inst_cell_71_125 ( BL125, BLN125, WL71);
sram_cell_6t_3 inst_cell_71_124 ( BL124, BLN124, WL71);
sram_cell_6t_3 inst_cell_71_123 ( BL123, BLN123, WL71);
sram_cell_6t_3 inst_cell_71_122 ( BL122, BLN122, WL71);
sram_cell_6t_3 inst_cell_71_121 ( BL121, BLN121, WL71);
sram_cell_6t_3 inst_cell_71_120 ( BL120, BLN120, WL71);
sram_cell_6t_3 inst_cell_71_119 ( BL119, BLN119, WL71);
sram_cell_6t_3 inst_cell_71_118 ( BL118, BLN118, WL71);
sram_cell_6t_3 inst_cell_71_117 ( BL117, BLN117, WL71);
sram_cell_6t_3 inst_cell_71_116 ( BL116, BLN116, WL71);
sram_cell_6t_3 inst_cell_71_115 ( BL115, BLN115, WL71);
sram_cell_6t_3 inst_cell_71_114 ( BL114, BLN114, WL71);
sram_cell_6t_3 inst_cell_71_113 ( BL113, BLN113, WL71);
sram_cell_6t_3 inst_cell_71_112 ( BL112, BLN112, WL71);
sram_cell_6t_3 inst_cell_71_111 ( BL111, BLN111, WL71);
sram_cell_6t_3 inst_cell_71_110 ( BL110, BLN110, WL71);
sram_cell_6t_3 inst_cell_71_109 ( BL109, BLN109, WL71);
sram_cell_6t_3 inst_cell_71_108 ( BL108, BLN108, WL71);
sram_cell_6t_3 inst_cell_71_107 ( BL107, BLN107, WL71);
sram_cell_6t_3 inst_cell_71_106 ( BL106, BLN106, WL71);
sram_cell_6t_3 inst_cell_71_105 ( BL105, BLN105, WL71);
sram_cell_6t_3 inst_cell_71_104 ( BL104, BLN104, WL71);
sram_cell_6t_3 inst_cell_71_103 ( BL103, BLN103, WL71);
sram_cell_6t_3 inst_cell_71_102 ( BL102, BLN102, WL71);
sram_cell_6t_3 inst_cell_71_101 ( BL101, BLN101, WL71);
sram_cell_6t_3 inst_cell_71_100 ( BL100, BLN100, WL71);
sram_cell_6t_3 inst_cell_71_99 ( BL99, BLN99, WL71);
sram_cell_6t_3 inst_cell_71_98 ( BL98, BLN98, WL71);
sram_cell_6t_3 inst_cell_71_97 ( BL97, BLN97, WL71);
sram_cell_6t_3 inst_cell_71_96 ( BL96, BLN96, WL71);
sram_cell_6t_3 inst_cell_71_95 ( BL95, BLN95, WL71);
sram_cell_6t_3 inst_cell_71_94 ( BL94, BLN94, WL71);
sram_cell_6t_3 inst_cell_71_93 ( BL93, BLN93, WL71);
sram_cell_6t_3 inst_cell_71_92 ( BL92, BLN92, WL71);
sram_cell_6t_3 inst_cell_71_91 ( BL91, BLN91, WL71);
sram_cell_6t_3 inst_cell_71_90 ( BL90, BLN90, WL71);
sram_cell_6t_3 inst_cell_71_89 ( BL89, BLN89, WL71);
sram_cell_6t_3 inst_cell_71_88 ( BL88, BLN88, WL71);
sram_cell_6t_3 inst_cell_71_87 ( BL87, BLN87, WL71);
sram_cell_6t_3 inst_cell_71_86 ( BL86, BLN86, WL71);
sram_cell_6t_3 inst_cell_71_85 ( BL85, BLN85, WL71);
sram_cell_6t_3 inst_cell_71_84 ( BL84, BLN84, WL71);
sram_cell_6t_3 inst_cell_71_83 ( BL83, BLN83, WL71);
sram_cell_6t_3 inst_cell_71_82 ( BL82, BLN82, WL71);
sram_cell_6t_3 inst_cell_71_81 ( BL81, BLN81, WL71);
sram_cell_6t_3 inst_cell_71_80 ( BL80, BLN80, WL71);
sram_cell_6t_3 inst_cell_71_79 ( BL79, BLN79, WL71);
sram_cell_6t_3 inst_cell_71_78 ( BL78, BLN78, WL71);
sram_cell_6t_3 inst_cell_71_77 ( BL77, BLN77, WL71);
sram_cell_6t_3 inst_cell_71_76 ( BL76, BLN76, WL71);
sram_cell_6t_3 inst_cell_71_75 ( BL75, BLN75, WL71);
sram_cell_6t_3 inst_cell_71_74 ( BL74, BLN74, WL71);
sram_cell_6t_3 inst_cell_71_73 ( BL73, BLN73, WL71);
sram_cell_6t_3 inst_cell_71_72 ( BL72, BLN72, WL71);
sram_cell_6t_3 inst_cell_71_71 ( BL71, BLN71, WL71);
sram_cell_6t_3 inst_cell_71_70 ( BL70, BLN70, WL71);
sram_cell_6t_3 inst_cell_71_69 ( BL69, BLN69, WL71);
sram_cell_6t_3 inst_cell_71_68 ( BL68, BLN68, WL71);
sram_cell_6t_3 inst_cell_71_67 ( BL67, BLN67, WL71);
sram_cell_6t_3 inst_cell_71_66 ( BL66, BLN66, WL71);
sram_cell_6t_3 inst_cell_71_65 ( BL65, BLN65, WL71);
sram_cell_6t_3 inst_cell_71_64 ( BL64, BLN64, WL71);
sram_cell_6t_3 inst_cell_71_63 ( BL63, BLN63, WL71);
sram_cell_6t_3 inst_cell_71_62 ( BL62, BLN62, WL71);
sram_cell_6t_3 inst_cell_71_61 ( BL61, BLN61, WL71);
sram_cell_6t_3 inst_cell_71_60 ( BL60, BLN60, WL71);
sram_cell_6t_3 inst_cell_71_59 ( BL59, BLN59, WL71);
sram_cell_6t_3 inst_cell_71_58 ( BL58, BLN58, WL71);
sram_cell_6t_3 inst_cell_71_57 ( BL57, BLN57, WL71);
sram_cell_6t_3 inst_cell_71_56 ( BL56, BLN56, WL71);
sram_cell_6t_3 inst_cell_71_55 ( BL55, BLN55, WL71);
sram_cell_6t_3 inst_cell_71_54 ( BL54, BLN54, WL71);
sram_cell_6t_3 inst_cell_71_53 ( BL53, BLN53, WL71);
sram_cell_6t_3 inst_cell_71_52 ( BL52, BLN52, WL71);
sram_cell_6t_3 inst_cell_71_51 ( BL51, BLN51, WL71);
sram_cell_6t_3 inst_cell_71_50 ( BL50, BLN50, WL71);
sram_cell_6t_3 inst_cell_71_49 ( BL49, BLN49, WL71);
sram_cell_6t_3 inst_cell_71_48 ( BL48, BLN48, WL71);
sram_cell_6t_3 inst_cell_71_47 ( BL47, BLN47, WL71);
sram_cell_6t_3 inst_cell_71_46 ( BL46, BLN46, WL71);
sram_cell_6t_3 inst_cell_71_45 ( BL45, BLN45, WL71);
sram_cell_6t_3 inst_cell_71_44 ( BL44, BLN44, WL71);
sram_cell_6t_3 inst_cell_71_43 ( BL43, BLN43, WL71);
sram_cell_6t_3 inst_cell_71_42 ( BL42, BLN42, WL71);
sram_cell_6t_3 inst_cell_71_41 ( BL41, BLN41, WL71);
sram_cell_6t_3 inst_cell_71_40 ( BL40, BLN40, WL71);
sram_cell_6t_3 inst_cell_71_39 ( BL39, BLN39, WL71);
sram_cell_6t_3 inst_cell_71_38 ( BL38, BLN38, WL71);
sram_cell_6t_3 inst_cell_71_37 ( BL37, BLN37, WL71);
sram_cell_6t_3 inst_cell_71_36 ( BL36, BLN36, WL71);
sram_cell_6t_3 inst_cell_71_35 ( BL35, BLN35, WL71);
sram_cell_6t_3 inst_cell_71_34 ( BL34, BLN34, WL71);
sram_cell_6t_3 inst_cell_71_33 ( BL33, BLN33, WL71);
sram_cell_6t_3 inst_cell_71_32 ( BL32, BLN32, WL71);
sram_cell_6t_3 inst_cell_71_31 ( BL31, BLN31, WL71);
sram_cell_6t_3 inst_cell_71_30 ( BL30, BLN30, WL71);
sram_cell_6t_3 inst_cell_71_29 ( BL29, BLN29, WL71);
sram_cell_6t_3 inst_cell_71_28 ( BL28, BLN28, WL71);
sram_cell_6t_3 inst_cell_71_27 ( BL27, BLN27, WL71);
sram_cell_6t_3 inst_cell_71_26 ( BL26, BLN26, WL71);
sram_cell_6t_3 inst_cell_71_25 ( BL25, BLN25, WL71);
sram_cell_6t_3 inst_cell_71_24 ( BL24, BLN24, WL71);
sram_cell_6t_3 inst_cell_71_23 ( BL23, BLN23, WL71);
sram_cell_6t_3 inst_cell_71_22 ( BL22, BLN22, WL71);
sram_cell_6t_3 inst_cell_71_21 ( BL21, BLN21, WL71);
sram_cell_6t_3 inst_cell_71_20 ( BL20, BLN20, WL71);
sram_cell_6t_3 inst_cell_71_19 ( BL19, BLN19, WL71);
sram_cell_6t_3 inst_cell_71_18 ( BL18, BLN18, WL71);
sram_cell_6t_3 inst_cell_71_17 ( BL17, BLN17, WL71);
sram_cell_6t_3 inst_cell_71_16 ( BL16, BLN16, WL71);
sram_cell_6t_3 inst_cell_71_15 ( BL15, BLN15, WL71);
sram_cell_6t_3 inst_cell_71_14 ( BL14, BLN14, WL71);
sram_cell_6t_3 inst_cell_71_13 ( BL13, BLN13, WL71);
sram_cell_6t_3 inst_cell_71_12 ( BL12, BLN12, WL71);
sram_cell_6t_3 inst_cell_71_11 ( BL11, BLN11, WL71);
sram_cell_6t_3 inst_cell_71_10 ( BL10, BLN10, WL71);
sram_cell_6t_3 inst_cell_71_9 ( BL9, BLN9, WL71);
sram_cell_6t_3 inst_cell_71_8 ( BL8, BLN8, WL71);
sram_cell_6t_3 inst_cell_71_7 ( BL7, BLN7, WL71);
sram_cell_6t_3 inst_cell_71_6 ( BL6, BLN6, WL71);
sram_cell_6t_3 inst_cell_71_5 ( BL5, BLN5, WL71);
sram_cell_6t_3 inst_cell_71_4 ( BL4, BLN4, WL71);
sram_cell_6t_3 inst_cell_71_3 ( BL3, BLN3, WL71);
sram_cell_6t_3 inst_cell_71_2 ( BL2, BLN2, WL71);
sram_cell_6t_3 inst_cell_71_1 ( BL1, BLN1, WL71);
sram_cell_6t_3 inst_cell_71_0 ( BL0, BLN0, WL71);
sram_cell_6t_3 inst_cell_70_127 ( BL127, BLN127, WL70);
sram_cell_6t_3 inst_cell_70_126 ( BL126, BLN126, WL70);
sram_cell_6t_3 inst_cell_70_125 ( BL125, BLN125, WL70);
sram_cell_6t_3 inst_cell_70_124 ( BL124, BLN124, WL70);
sram_cell_6t_3 inst_cell_70_123 ( BL123, BLN123, WL70);
sram_cell_6t_3 inst_cell_70_122 ( BL122, BLN122, WL70);
sram_cell_6t_3 inst_cell_70_121 ( BL121, BLN121, WL70);
sram_cell_6t_3 inst_cell_70_120 ( BL120, BLN120, WL70);
sram_cell_6t_3 inst_cell_70_119 ( BL119, BLN119, WL70);
sram_cell_6t_3 inst_cell_70_118 ( BL118, BLN118, WL70);
sram_cell_6t_3 inst_cell_70_117 ( BL117, BLN117, WL70);
sram_cell_6t_3 inst_cell_70_116 ( BL116, BLN116, WL70);
sram_cell_6t_3 inst_cell_70_115 ( BL115, BLN115, WL70);
sram_cell_6t_3 inst_cell_70_114 ( BL114, BLN114, WL70);
sram_cell_6t_3 inst_cell_70_113 ( BL113, BLN113, WL70);
sram_cell_6t_3 inst_cell_70_112 ( BL112, BLN112, WL70);
sram_cell_6t_3 inst_cell_70_111 ( BL111, BLN111, WL70);
sram_cell_6t_3 inst_cell_70_110 ( BL110, BLN110, WL70);
sram_cell_6t_3 inst_cell_70_109 ( BL109, BLN109, WL70);
sram_cell_6t_3 inst_cell_70_108 ( BL108, BLN108, WL70);
sram_cell_6t_3 inst_cell_70_107 ( BL107, BLN107, WL70);
sram_cell_6t_3 inst_cell_70_106 ( BL106, BLN106, WL70);
sram_cell_6t_3 inst_cell_70_105 ( BL105, BLN105, WL70);
sram_cell_6t_3 inst_cell_70_104 ( BL104, BLN104, WL70);
sram_cell_6t_3 inst_cell_70_103 ( BL103, BLN103, WL70);
sram_cell_6t_3 inst_cell_70_102 ( BL102, BLN102, WL70);
sram_cell_6t_3 inst_cell_70_101 ( BL101, BLN101, WL70);
sram_cell_6t_3 inst_cell_70_100 ( BL100, BLN100, WL70);
sram_cell_6t_3 inst_cell_70_99 ( BL99, BLN99, WL70);
sram_cell_6t_3 inst_cell_70_98 ( BL98, BLN98, WL70);
sram_cell_6t_3 inst_cell_70_97 ( BL97, BLN97, WL70);
sram_cell_6t_3 inst_cell_70_96 ( BL96, BLN96, WL70);
sram_cell_6t_3 inst_cell_70_95 ( BL95, BLN95, WL70);
sram_cell_6t_3 inst_cell_70_94 ( BL94, BLN94, WL70);
sram_cell_6t_3 inst_cell_70_93 ( BL93, BLN93, WL70);
sram_cell_6t_3 inst_cell_70_92 ( BL92, BLN92, WL70);
sram_cell_6t_3 inst_cell_70_91 ( BL91, BLN91, WL70);
sram_cell_6t_3 inst_cell_70_90 ( BL90, BLN90, WL70);
sram_cell_6t_3 inst_cell_70_89 ( BL89, BLN89, WL70);
sram_cell_6t_3 inst_cell_70_88 ( BL88, BLN88, WL70);
sram_cell_6t_3 inst_cell_70_87 ( BL87, BLN87, WL70);
sram_cell_6t_3 inst_cell_70_86 ( BL86, BLN86, WL70);
sram_cell_6t_3 inst_cell_70_85 ( BL85, BLN85, WL70);
sram_cell_6t_3 inst_cell_70_84 ( BL84, BLN84, WL70);
sram_cell_6t_3 inst_cell_70_83 ( BL83, BLN83, WL70);
sram_cell_6t_3 inst_cell_70_82 ( BL82, BLN82, WL70);
sram_cell_6t_3 inst_cell_70_81 ( BL81, BLN81, WL70);
sram_cell_6t_3 inst_cell_70_80 ( BL80, BLN80, WL70);
sram_cell_6t_3 inst_cell_70_79 ( BL79, BLN79, WL70);
sram_cell_6t_3 inst_cell_70_78 ( BL78, BLN78, WL70);
sram_cell_6t_3 inst_cell_70_77 ( BL77, BLN77, WL70);
sram_cell_6t_3 inst_cell_70_76 ( BL76, BLN76, WL70);
sram_cell_6t_3 inst_cell_70_75 ( BL75, BLN75, WL70);
sram_cell_6t_3 inst_cell_70_74 ( BL74, BLN74, WL70);
sram_cell_6t_3 inst_cell_70_73 ( BL73, BLN73, WL70);
sram_cell_6t_3 inst_cell_70_72 ( BL72, BLN72, WL70);
sram_cell_6t_3 inst_cell_70_71 ( BL71, BLN71, WL70);
sram_cell_6t_3 inst_cell_70_70 ( BL70, BLN70, WL70);
sram_cell_6t_3 inst_cell_70_69 ( BL69, BLN69, WL70);
sram_cell_6t_3 inst_cell_70_68 ( BL68, BLN68, WL70);
sram_cell_6t_3 inst_cell_70_67 ( BL67, BLN67, WL70);
sram_cell_6t_3 inst_cell_70_66 ( BL66, BLN66, WL70);
sram_cell_6t_3 inst_cell_70_65 ( BL65, BLN65, WL70);
sram_cell_6t_3 inst_cell_70_64 ( BL64, BLN64, WL70);
sram_cell_6t_3 inst_cell_70_63 ( BL63, BLN63, WL70);
sram_cell_6t_3 inst_cell_70_62 ( BL62, BLN62, WL70);
sram_cell_6t_3 inst_cell_70_61 ( BL61, BLN61, WL70);
sram_cell_6t_3 inst_cell_70_60 ( BL60, BLN60, WL70);
sram_cell_6t_3 inst_cell_70_59 ( BL59, BLN59, WL70);
sram_cell_6t_3 inst_cell_70_58 ( BL58, BLN58, WL70);
sram_cell_6t_3 inst_cell_70_57 ( BL57, BLN57, WL70);
sram_cell_6t_3 inst_cell_70_56 ( BL56, BLN56, WL70);
sram_cell_6t_3 inst_cell_70_55 ( BL55, BLN55, WL70);
sram_cell_6t_3 inst_cell_70_54 ( BL54, BLN54, WL70);
sram_cell_6t_3 inst_cell_70_53 ( BL53, BLN53, WL70);
sram_cell_6t_3 inst_cell_70_52 ( BL52, BLN52, WL70);
sram_cell_6t_3 inst_cell_70_51 ( BL51, BLN51, WL70);
sram_cell_6t_3 inst_cell_70_50 ( BL50, BLN50, WL70);
sram_cell_6t_3 inst_cell_70_49 ( BL49, BLN49, WL70);
sram_cell_6t_3 inst_cell_70_48 ( BL48, BLN48, WL70);
sram_cell_6t_3 inst_cell_70_47 ( BL47, BLN47, WL70);
sram_cell_6t_3 inst_cell_70_46 ( BL46, BLN46, WL70);
sram_cell_6t_3 inst_cell_70_45 ( BL45, BLN45, WL70);
sram_cell_6t_3 inst_cell_70_44 ( BL44, BLN44, WL70);
sram_cell_6t_3 inst_cell_70_43 ( BL43, BLN43, WL70);
sram_cell_6t_3 inst_cell_70_42 ( BL42, BLN42, WL70);
sram_cell_6t_3 inst_cell_70_41 ( BL41, BLN41, WL70);
sram_cell_6t_3 inst_cell_70_40 ( BL40, BLN40, WL70);
sram_cell_6t_3 inst_cell_70_39 ( BL39, BLN39, WL70);
sram_cell_6t_3 inst_cell_70_38 ( BL38, BLN38, WL70);
sram_cell_6t_3 inst_cell_70_37 ( BL37, BLN37, WL70);
sram_cell_6t_3 inst_cell_70_36 ( BL36, BLN36, WL70);
sram_cell_6t_3 inst_cell_70_35 ( BL35, BLN35, WL70);
sram_cell_6t_3 inst_cell_70_34 ( BL34, BLN34, WL70);
sram_cell_6t_3 inst_cell_70_33 ( BL33, BLN33, WL70);
sram_cell_6t_3 inst_cell_70_32 ( BL32, BLN32, WL70);
sram_cell_6t_3 inst_cell_70_31 ( BL31, BLN31, WL70);
sram_cell_6t_3 inst_cell_70_30 ( BL30, BLN30, WL70);
sram_cell_6t_3 inst_cell_70_29 ( BL29, BLN29, WL70);
sram_cell_6t_3 inst_cell_70_28 ( BL28, BLN28, WL70);
sram_cell_6t_3 inst_cell_70_27 ( BL27, BLN27, WL70);
sram_cell_6t_3 inst_cell_70_26 ( BL26, BLN26, WL70);
sram_cell_6t_3 inst_cell_70_25 ( BL25, BLN25, WL70);
sram_cell_6t_3 inst_cell_70_24 ( BL24, BLN24, WL70);
sram_cell_6t_3 inst_cell_70_23 ( BL23, BLN23, WL70);
sram_cell_6t_3 inst_cell_70_22 ( BL22, BLN22, WL70);
sram_cell_6t_3 inst_cell_70_21 ( BL21, BLN21, WL70);
sram_cell_6t_3 inst_cell_70_20 ( BL20, BLN20, WL70);
sram_cell_6t_3 inst_cell_70_19 ( BL19, BLN19, WL70);
sram_cell_6t_3 inst_cell_70_18 ( BL18, BLN18, WL70);
sram_cell_6t_3 inst_cell_70_17 ( BL17, BLN17, WL70);
sram_cell_6t_3 inst_cell_70_16 ( BL16, BLN16, WL70);
sram_cell_6t_3 inst_cell_70_15 ( BL15, BLN15, WL70);
sram_cell_6t_3 inst_cell_70_14 ( BL14, BLN14, WL70);
sram_cell_6t_3 inst_cell_70_13 ( BL13, BLN13, WL70);
sram_cell_6t_3 inst_cell_70_12 ( BL12, BLN12, WL70);
sram_cell_6t_3 inst_cell_70_11 ( BL11, BLN11, WL70);
sram_cell_6t_3 inst_cell_70_10 ( BL10, BLN10, WL70);
sram_cell_6t_3 inst_cell_70_9 ( BL9, BLN9, WL70);
sram_cell_6t_3 inst_cell_70_8 ( BL8, BLN8, WL70);
sram_cell_6t_3 inst_cell_70_7 ( BL7, BLN7, WL70);
sram_cell_6t_3 inst_cell_70_6 ( BL6, BLN6, WL70);
sram_cell_6t_3 inst_cell_70_5 ( BL5, BLN5, WL70);
sram_cell_6t_3 inst_cell_70_4 ( BL4, BLN4, WL70);
sram_cell_6t_3 inst_cell_70_3 ( BL3, BLN3, WL70);
sram_cell_6t_3 inst_cell_70_2 ( BL2, BLN2, WL70);
sram_cell_6t_3 inst_cell_70_1 ( BL1, BLN1, WL70);
sram_cell_6t_3 inst_cell_70_0 ( BL0, BLN0, WL70);
sram_cell_6t_3 inst_cell_69_127 ( BL127, BLN127, WL69);
sram_cell_6t_3 inst_cell_69_126 ( BL126, BLN126, WL69);
sram_cell_6t_3 inst_cell_69_125 ( BL125, BLN125, WL69);
sram_cell_6t_3 inst_cell_69_124 ( BL124, BLN124, WL69);
sram_cell_6t_3 inst_cell_69_123 ( BL123, BLN123, WL69);
sram_cell_6t_3 inst_cell_69_122 ( BL122, BLN122, WL69);
sram_cell_6t_3 inst_cell_69_121 ( BL121, BLN121, WL69);
sram_cell_6t_3 inst_cell_69_120 ( BL120, BLN120, WL69);
sram_cell_6t_3 inst_cell_69_119 ( BL119, BLN119, WL69);
sram_cell_6t_3 inst_cell_69_118 ( BL118, BLN118, WL69);
sram_cell_6t_3 inst_cell_69_117 ( BL117, BLN117, WL69);
sram_cell_6t_3 inst_cell_69_116 ( BL116, BLN116, WL69);
sram_cell_6t_3 inst_cell_69_115 ( BL115, BLN115, WL69);
sram_cell_6t_3 inst_cell_69_114 ( BL114, BLN114, WL69);
sram_cell_6t_3 inst_cell_69_113 ( BL113, BLN113, WL69);
sram_cell_6t_3 inst_cell_69_112 ( BL112, BLN112, WL69);
sram_cell_6t_3 inst_cell_69_111 ( BL111, BLN111, WL69);
sram_cell_6t_3 inst_cell_69_110 ( BL110, BLN110, WL69);
sram_cell_6t_3 inst_cell_69_109 ( BL109, BLN109, WL69);
sram_cell_6t_3 inst_cell_69_108 ( BL108, BLN108, WL69);
sram_cell_6t_3 inst_cell_69_107 ( BL107, BLN107, WL69);
sram_cell_6t_3 inst_cell_69_106 ( BL106, BLN106, WL69);
sram_cell_6t_3 inst_cell_69_105 ( BL105, BLN105, WL69);
sram_cell_6t_3 inst_cell_69_104 ( BL104, BLN104, WL69);
sram_cell_6t_3 inst_cell_69_103 ( BL103, BLN103, WL69);
sram_cell_6t_3 inst_cell_69_102 ( BL102, BLN102, WL69);
sram_cell_6t_3 inst_cell_69_101 ( BL101, BLN101, WL69);
sram_cell_6t_3 inst_cell_69_100 ( BL100, BLN100, WL69);
sram_cell_6t_3 inst_cell_69_99 ( BL99, BLN99, WL69);
sram_cell_6t_3 inst_cell_69_98 ( BL98, BLN98, WL69);
sram_cell_6t_3 inst_cell_69_97 ( BL97, BLN97, WL69);
sram_cell_6t_3 inst_cell_69_96 ( BL96, BLN96, WL69);
sram_cell_6t_3 inst_cell_69_95 ( BL95, BLN95, WL69);
sram_cell_6t_3 inst_cell_69_94 ( BL94, BLN94, WL69);
sram_cell_6t_3 inst_cell_69_93 ( BL93, BLN93, WL69);
sram_cell_6t_3 inst_cell_69_92 ( BL92, BLN92, WL69);
sram_cell_6t_3 inst_cell_69_91 ( BL91, BLN91, WL69);
sram_cell_6t_3 inst_cell_69_90 ( BL90, BLN90, WL69);
sram_cell_6t_3 inst_cell_69_89 ( BL89, BLN89, WL69);
sram_cell_6t_3 inst_cell_69_88 ( BL88, BLN88, WL69);
sram_cell_6t_3 inst_cell_69_87 ( BL87, BLN87, WL69);
sram_cell_6t_3 inst_cell_69_86 ( BL86, BLN86, WL69);
sram_cell_6t_3 inst_cell_69_85 ( BL85, BLN85, WL69);
sram_cell_6t_3 inst_cell_69_84 ( BL84, BLN84, WL69);
sram_cell_6t_3 inst_cell_69_83 ( BL83, BLN83, WL69);
sram_cell_6t_3 inst_cell_69_82 ( BL82, BLN82, WL69);
sram_cell_6t_3 inst_cell_69_81 ( BL81, BLN81, WL69);
sram_cell_6t_3 inst_cell_69_80 ( BL80, BLN80, WL69);
sram_cell_6t_3 inst_cell_69_79 ( BL79, BLN79, WL69);
sram_cell_6t_3 inst_cell_69_78 ( BL78, BLN78, WL69);
sram_cell_6t_3 inst_cell_69_77 ( BL77, BLN77, WL69);
sram_cell_6t_3 inst_cell_69_76 ( BL76, BLN76, WL69);
sram_cell_6t_3 inst_cell_69_75 ( BL75, BLN75, WL69);
sram_cell_6t_3 inst_cell_69_74 ( BL74, BLN74, WL69);
sram_cell_6t_3 inst_cell_69_73 ( BL73, BLN73, WL69);
sram_cell_6t_3 inst_cell_69_72 ( BL72, BLN72, WL69);
sram_cell_6t_3 inst_cell_69_71 ( BL71, BLN71, WL69);
sram_cell_6t_3 inst_cell_69_70 ( BL70, BLN70, WL69);
sram_cell_6t_3 inst_cell_69_69 ( BL69, BLN69, WL69);
sram_cell_6t_3 inst_cell_69_68 ( BL68, BLN68, WL69);
sram_cell_6t_3 inst_cell_69_67 ( BL67, BLN67, WL69);
sram_cell_6t_3 inst_cell_69_66 ( BL66, BLN66, WL69);
sram_cell_6t_3 inst_cell_69_65 ( BL65, BLN65, WL69);
sram_cell_6t_3 inst_cell_69_64 ( BL64, BLN64, WL69);
sram_cell_6t_3 inst_cell_69_63 ( BL63, BLN63, WL69);
sram_cell_6t_3 inst_cell_69_62 ( BL62, BLN62, WL69);
sram_cell_6t_3 inst_cell_69_61 ( BL61, BLN61, WL69);
sram_cell_6t_3 inst_cell_69_60 ( BL60, BLN60, WL69);
sram_cell_6t_3 inst_cell_69_59 ( BL59, BLN59, WL69);
sram_cell_6t_3 inst_cell_69_58 ( BL58, BLN58, WL69);
sram_cell_6t_3 inst_cell_69_57 ( BL57, BLN57, WL69);
sram_cell_6t_3 inst_cell_69_56 ( BL56, BLN56, WL69);
sram_cell_6t_3 inst_cell_69_55 ( BL55, BLN55, WL69);
sram_cell_6t_3 inst_cell_69_54 ( BL54, BLN54, WL69);
sram_cell_6t_3 inst_cell_69_53 ( BL53, BLN53, WL69);
sram_cell_6t_3 inst_cell_69_52 ( BL52, BLN52, WL69);
sram_cell_6t_3 inst_cell_69_51 ( BL51, BLN51, WL69);
sram_cell_6t_3 inst_cell_69_50 ( BL50, BLN50, WL69);
sram_cell_6t_3 inst_cell_69_49 ( BL49, BLN49, WL69);
sram_cell_6t_3 inst_cell_69_48 ( BL48, BLN48, WL69);
sram_cell_6t_3 inst_cell_69_47 ( BL47, BLN47, WL69);
sram_cell_6t_3 inst_cell_69_46 ( BL46, BLN46, WL69);
sram_cell_6t_3 inst_cell_69_45 ( BL45, BLN45, WL69);
sram_cell_6t_3 inst_cell_69_44 ( BL44, BLN44, WL69);
sram_cell_6t_3 inst_cell_69_43 ( BL43, BLN43, WL69);
sram_cell_6t_3 inst_cell_69_42 ( BL42, BLN42, WL69);
sram_cell_6t_3 inst_cell_69_41 ( BL41, BLN41, WL69);
sram_cell_6t_3 inst_cell_69_40 ( BL40, BLN40, WL69);
sram_cell_6t_3 inst_cell_69_39 ( BL39, BLN39, WL69);
sram_cell_6t_3 inst_cell_69_38 ( BL38, BLN38, WL69);
sram_cell_6t_3 inst_cell_69_37 ( BL37, BLN37, WL69);
sram_cell_6t_3 inst_cell_69_36 ( BL36, BLN36, WL69);
sram_cell_6t_3 inst_cell_69_35 ( BL35, BLN35, WL69);
sram_cell_6t_3 inst_cell_69_34 ( BL34, BLN34, WL69);
sram_cell_6t_3 inst_cell_69_33 ( BL33, BLN33, WL69);
sram_cell_6t_3 inst_cell_69_32 ( BL32, BLN32, WL69);
sram_cell_6t_3 inst_cell_69_31 ( BL31, BLN31, WL69);
sram_cell_6t_3 inst_cell_69_30 ( BL30, BLN30, WL69);
sram_cell_6t_3 inst_cell_69_29 ( BL29, BLN29, WL69);
sram_cell_6t_3 inst_cell_69_28 ( BL28, BLN28, WL69);
sram_cell_6t_3 inst_cell_69_27 ( BL27, BLN27, WL69);
sram_cell_6t_3 inst_cell_69_26 ( BL26, BLN26, WL69);
sram_cell_6t_3 inst_cell_69_25 ( BL25, BLN25, WL69);
sram_cell_6t_3 inst_cell_69_24 ( BL24, BLN24, WL69);
sram_cell_6t_3 inst_cell_69_23 ( BL23, BLN23, WL69);
sram_cell_6t_3 inst_cell_69_22 ( BL22, BLN22, WL69);
sram_cell_6t_3 inst_cell_69_21 ( BL21, BLN21, WL69);
sram_cell_6t_3 inst_cell_69_20 ( BL20, BLN20, WL69);
sram_cell_6t_3 inst_cell_69_19 ( BL19, BLN19, WL69);
sram_cell_6t_3 inst_cell_69_18 ( BL18, BLN18, WL69);
sram_cell_6t_3 inst_cell_69_17 ( BL17, BLN17, WL69);
sram_cell_6t_3 inst_cell_69_16 ( BL16, BLN16, WL69);
sram_cell_6t_3 inst_cell_69_15 ( BL15, BLN15, WL69);
sram_cell_6t_3 inst_cell_69_14 ( BL14, BLN14, WL69);
sram_cell_6t_3 inst_cell_69_13 ( BL13, BLN13, WL69);
sram_cell_6t_3 inst_cell_69_12 ( BL12, BLN12, WL69);
sram_cell_6t_3 inst_cell_69_11 ( BL11, BLN11, WL69);
sram_cell_6t_3 inst_cell_69_10 ( BL10, BLN10, WL69);
sram_cell_6t_3 inst_cell_69_9 ( BL9, BLN9, WL69);
sram_cell_6t_3 inst_cell_69_8 ( BL8, BLN8, WL69);
sram_cell_6t_3 inst_cell_69_7 ( BL7, BLN7, WL69);
sram_cell_6t_3 inst_cell_69_6 ( BL6, BLN6, WL69);
sram_cell_6t_3 inst_cell_69_5 ( BL5, BLN5, WL69);
sram_cell_6t_3 inst_cell_69_4 ( BL4, BLN4, WL69);
sram_cell_6t_3 inst_cell_69_3 ( BL3, BLN3, WL69);
sram_cell_6t_3 inst_cell_69_2 ( BL2, BLN2, WL69);
sram_cell_6t_3 inst_cell_69_1 ( BL1, BLN1, WL69);
sram_cell_6t_3 inst_cell_69_0 ( BL0, BLN0, WL69);
sram_cell_6t_3 inst_cell_68_127 ( BL127, BLN127, WL68);
sram_cell_6t_3 inst_cell_68_126 ( BL126, BLN126, WL68);
sram_cell_6t_3 inst_cell_68_125 ( BL125, BLN125, WL68);
sram_cell_6t_3 inst_cell_68_124 ( BL124, BLN124, WL68);
sram_cell_6t_3 inst_cell_68_123 ( BL123, BLN123, WL68);
sram_cell_6t_3 inst_cell_68_122 ( BL122, BLN122, WL68);
sram_cell_6t_3 inst_cell_68_121 ( BL121, BLN121, WL68);
sram_cell_6t_3 inst_cell_68_120 ( BL120, BLN120, WL68);
sram_cell_6t_3 inst_cell_68_119 ( BL119, BLN119, WL68);
sram_cell_6t_3 inst_cell_68_118 ( BL118, BLN118, WL68);
sram_cell_6t_3 inst_cell_68_117 ( BL117, BLN117, WL68);
sram_cell_6t_3 inst_cell_68_116 ( BL116, BLN116, WL68);
sram_cell_6t_3 inst_cell_68_115 ( BL115, BLN115, WL68);
sram_cell_6t_3 inst_cell_68_114 ( BL114, BLN114, WL68);
sram_cell_6t_3 inst_cell_68_113 ( BL113, BLN113, WL68);
sram_cell_6t_3 inst_cell_68_112 ( BL112, BLN112, WL68);
sram_cell_6t_3 inst_cell_68_111 ( BL111, BLN111, WL68);
sram_cell_6t_3 inst_cell_68_110 ( BL110, BLN110, WL68);
sram_cell_6t_3 inst_cell_68_109 ( BL109, BLN109, WL68);
sram_cell_6t_3 inst_cell_68_108 ( BL108, BLN108, WL68);
sram_cell_6t_3 inst_cell_68_107 ( BL107, BLN107, WL68);
sram_cell_6t_3 inst_cell_68_106 ( BL106, BLN106, WL68);
sram_cell_6t_3 inst_cell_68_105 ( BL105, BLN105, WL68);
sram_cell_6t_3 inst_cell_68_104 ( BL104, BLN104, WL68);
sram_cell_6t_3 inst_cell_68_103 ( BL103, BLN103, WL68);
sram_cell_6t_3 inst_cell_68_102 ( BL102, BLN102, WL68);
sram_cell_6t_3 inst_cell_68_101 ( BL101, BLN101, WL68);
sram_cell_6t_3 inst_cell_68_100 ( BL100, BLN100, WL68);
sram_cell_6t_3 inst_cell_68_99 ( BL99, BLN99, WL68);
sram_cell_6t_3 inst_cell_68_98 ( BL98, BLN98, WL68);
sram_cell_6t_3 inst_cell_68_97 ( BL97, BLN97, WL68);
sram_cell_6t_3 inst_cell_68_96 ( BL96, BLN96, WL68);
sram_cell_6t_3 inst_cell_68_95 ( BL95, BLN95, WL68);
sram_cell_6t_3 inst_cell_68_94 ( BL94, BLN94, WL68);
sram_cell_6t_3 inst_cell_68_93 ( BL93, BLN93, WL68);
sram_cell_6t_3 inst_cell_68_92 ( BL92, BLN92, WL68);
sram_cell_6t_3 inst_cell_68_91 ( BL91, BLN91, WL68);
sram_cell_6t_3 inst_cell_68_90 ( BL90, BLN90, WL68);
sram_cell_6t_3 inst_cell_68_89 ( BL89, BLN89, WL68);
sram_cell_6t_3 inst_cell_68_88 ( BL88, BLN88, WL68);
sram_cell_6t_3 inst_cell_68_87 ( BL87, BLN87, WL68);
sram_cell_6t_3 inst_cell_68_86 ( BL86, BLN86, WL68);
sram_cell_6t_3 inst_cell_68_85 ( BL85, BLN85, WL68);
sram_cell_6t_3 inst_cell_68_84 ( BL84, BLN84, WL68);
sram_cell_6t_3 inst_cell_68_83 ( BL83, BLN83, WL68);
sram_cell_6t_3 inst_cell_68_82 ( BL82, BLN82, WL68);
sram_cell_6t_3 inst_cell_68_81 ( BL81, BLN81, WL68);
sram_cell_6t_3 inst_cell_68_80 ( BL80, BLN80, WL68);
sram_cell_6t_3 inst_cell_68_79 ( BL79, BLN79, WL68);
sram_cell_6t_3 inst_cell_68_78 ( BL78, BLN78, WL68);
sram_cell_6t_3 inst_cell_68_77 ( BL77, BLN77, WL68);
sram_cell_6t_3 inst_cell_68_76 ( BL76, BLN76, WL68);
sram_cell_6t_3 inst_cell_68_75 ( BL75, BLN75, WL68);
sram_cell_6t_3 inst_cell_68_74 ( BL74, BLN74, WL68);
sram_cell_6t_3 inst_cell_68_73 ( BL73, BLN73, WL68);
sram_cell_6t_3 inst_cell_68_72 ( BL72, BLN72, WL68);
sram_cell_6t_3 inst_cell_68_71 ( BL71, BLN71, WL68);
sram_cell_6t_3 inst_cell_68_70 ( BL70, BLN70, WL68);
sram_cell_6t_3 inst_cell_68_69 ( BL69, BLN69, WL68);
sram_cell_6t_3 inst_cell_68_68 ( BL68, BLN68, WL68);
sram_cell_6t_3 inst_cell_68_67 ( BL67, BLN67, WL68);
sram_cell_6t_3 inst_cell_68_66 ( BL66, BLN66, WL68);
sram_cell_6t_3 inst_cell_68_65 ( BL65, BLN65, WL68);
sram_cell_6t_3 inst_cell_68_64 ( BL64, BLN64, WL68);
sram_cell_6t_3 inst_cell_68_63 ( BL63, BLN63, WL68);
sram_cell_6t_3 inst_cell_68_62 ( BL62, BLN62, WL68);
sram_cell_6t_3 inst_cell_68_61 ( BL61, BLN61, WL68);
sram_cell_6t_3 inst_cell_68_60 ( BL60, BLN60, WL68);
sram_cell_6t_3 inst_cell_68_59 ( BL59, BLN59, WL68);
sram_cell_6t_3 inst_cell_68_58 ( BL58, BLN58, WL68);
sram_cell_6t_3 inst_cell_68_57 ( BL57, BLN57, WL68);
sram_cell_6t_3 inst_cell_68_56 ( BL56, BLN56, WL68);
sram_cell_6t_3 inst_cell_68_55 ( BL55, BLN55, WL68);
sram_cell_6t_3 inst_cell_68_54 ( BL54, BLN54, WL68);
sram_cell_6t_3 inst_cell_68_53 ( BL53, BLN53, WL68);
sram_cell_6t_3 inst_cell_68_52 ( BL52, BLN52, WL68);
sram_cell_6t_3 inst_cell_68_51 ( BL51, BLN51, WL68);
sram_cell_6t_3 inst_cell_68_50 ( BL50, BLN50, WL68);
sram_cell_6t_3 inst_cell_68_49 ( BL49, BLN49, WL68);
sram_cell_6t_3 inst_cell_68_48 ( BL48, BLN48, WL68);
sram_cell_6t_3 inst_cell_68_47 ( BL47, BLN47, WL68);
sram_cell_6t_3 inst_cell_68_46 ( BL46, BLN46, WL68);
sram_cell_6t_3 inst_cell_68_45 ( BL45, BLN45, WL68);
sram_cell_6t_3 inst_cell_68_44 ( BL44, BLN44, WL68);
sram_cell_6t_3 inst_cell_68_43 ( BL43, BLN43, WL68);
sram_cell_6t_3 inst_cell_68_42 ( BL42, BLN42, WL68);
sram_cell_6t_3 inst_cell_68_41 ( BL41, BLN41, WL68);
sram_cell_6t_3 inst_cell_68_40 ( BL40, BLN40, WL68);
sram_cell_6t_3 inst_cell_68_39 ( BL39, BLN39, WL68);
sram_cell_6t_3 inst_cell_68_38 ( BL38, BLN38, WL68);
sram_cell_6t_3 inst_cell_68_37 ( BL37, BLN37, WL68);
sram_cell_6t_3 inst_cell_68_36 ( BL36, BLN36, WL68);
sram_cell_6t_3 inst_cell_68_35 ( BL35, BLN35, WL68);
sram_cell_6t_3 inst_cell_68_34 ( BL34, BLN34, WL68);
sram_cell_6t_3 inst_cell_68_33 ( BL33, BLN33, WL68);
sram_cell_6t_3 inst_cell_68_32 ( BL32, BLN32, WL68);
sram_cell_6t_3 inst_cell_68_31 ( BL31, BLN31, WL68);
sram_cell_6t_3 inst_cell_68_30 ( BL30, BLN30, WL68);
sram_cell_6t_3 inst_cell_68_29 ( BL29, BLN29, WL68);
sram_cell_6t_3 inst_cell_68_28 ( BL28, BLN28, WL68);
sram_cell_6t_3 inst_cell_68_27 ( BL27, BLN27, WL68);
sram_cell_6t_3 inst_cell_68_26 ( BL26, BLN26, WL68);
sram_cell_6t_3 inst_cell_68_25 ( BL25, BLN25, WL68);
sram_cell_6t_3 inst_cell_68_24 ( BL24, BLN24, WL68);
sram_cell_6t_3 inst_cell_68_23 ( BL23, BLN23, WL68);
sram_cell_6t_3 inst_cell_68_22 ( BL22, BLN22, WL68);
sram_cell_6t_3 inst_cell_68_21 ( BL21, BLN21, WL68);
sram_cell_6t_3 inst_cell_68_20 ( BL20, BLN20, WL68);
sram_cell_6t_3 inst_cell_68_19 ( BL19, BLN19, WL68);
sram_cell_6t_3 inst_cell_68_18 ( BL18, BLN18, WL68);
sram_cell_6t_3 inst_cell_68_17 ( BL17, BLN17, WL68);
sram_cell_6t_3 inst_cell_68_16 ( BL16, BLN16, WL68);
sram_cell_6t_3 inst_cell_68_15 ( BL15, BLN15, WL68);
sram_cell_6t_3 inst_cell_68_14 ( BL14, BLN14, WL68);
sram_cell_6t_3 inst_cell_68_13 ( BL13, BLN13, WL68);
sram_cell_6t_3 inst_cell_68_12 ( BL12, BLN12, WL68);
sram_cell_6t_3 inst_cell_68_11 ( BL11, BLN11, WL68);
sram_cell_6t_3 inst_cell_68_10 ( BL10, BLN10, WL68);
sram_cell_6t_3 inst_cell_68_9 ( BL9, BLN9, WL68);
sram_cell_6t_3 inst_cell_68_8 ( BL8, BLN8, WL68);
sram_cell_6t_3 inst_cell_68_7 ( BL7, BLN7, WL68);
sram_cell_6t_3 inst_cell_68_6 ( BL6, BLN6, WL68);
sram_cell_6t_3 inst_cell_68_5 ( BL5, BLN5, WL68);
sram_cell_6t_3 inst_cell_68_4 ( BL4, BLN4, WL68);
sram_cell_6t_3 inst_cell_68_3 ( BL3, BLN3, WL68);
sram_cell_6t_3 inst_cell_68_2 ( BL2, BLN2, WL68);
sram_cell_6t_3 inst_cell_68_1 ( BL1, BLN1, WL68);
sram_cell_6t_3 inst_cell_68_0 ( BL0, BLN0, WL68);
sram_cell_6t_3 inst_cell_67_127 ( BL127, BLN127, WL67);
sram_cell_6t_3 inst_cell_67_126 ( BL126, BLN126, WL67);
sram_cell_6t_3 inst_cell_67_125 ( BL125, BLN125, WL67);
sram_cell_6t_3 inst_cell_67_124 ( BL124, BLN124, WL67);
sram_cell_6t_3 inst_cell_67_123 ( BL123, BLN123, WL67);
sram_cell_6t_3 inst_cell_67_122 ( BL122, BLN122, WL67);
sram_cell_6t_3 inst_cell_67_121 ( BL121, BLN121, WL67);
sram_cell_6t_3 inst_cell_67_120 ( BL120, BLN120, WL67);
sram_cell_6t_3 inst_cell_67_119 ( BL119, BLN119, WL67);
sram_cell_6t_3 inst_cell_67_118 ( BL118, BLN118, WL67);
sram_cell_6t_3 inst_cell_67_117 ( BL117, BLN117, WL67);
sram_cell_6t_3 inst_cell_67_116 ( BL116, BLN116, WL67);
sram_cell_6t_3 inst_cell_67_115 ( BL115, BLN115, WL67);
sram_cell_6t_3 inst_cell_67_114 ( BL114, BLN114, WL67);
sram_cell_6t_3 inst_cell_67_113 ( BL113, BLN113, WL67);
sram_cell_6t_3 inst_cell_67_112 ( BL112, BLN112, WL67);
sram_cell_6t_3 inst_cell_67_111 ( BL111, BLN111, WL67);
sram_cell_6t_3 inst_cell_67_110 ( BL110, BLN110, WL67);
sram_cell_6t_3 inst_cell_67_109 ( BL109, BLN109, WL67);
sram_cell_6t_3 inst_cell_67_108 ( BL108, BLN108, WL67);
sram_cell_6t_3 inst_cell_67_107 ( BL107, BLN107, WL67);
sram_cell_6t_3 inst_cell_67_106 ( BL106, BLN106, WL67);
sram_cell_6t_3 inst_cell_67_105 ( BL105, BLN105, WL67);
sram_cell_6t_3 inst_cell_67_104 ( BL104, BLN104, WL67);
sram_cell_6t_3 inst_cell_67_103 ( BL103, BLN103, WL67);
sram_cell_6t_3 inst_cell_67_102 ( BL102, BLN102, WL67);
sram_cell_6t_3 inst_cell_67_101 ( BL101, BLN101, WL67);
sram_cell_6t_3 inst_cell_67_100 ( BL100, BLN100, WL67);
sram_cell_6t_3 inst_cell_67_99 ( BL99, BLN99, WL67);
sram_cell_6t_3 inst_cell_67_98 ( BL98, BLN98, WL67);
sram_cell_6t_3 inst_cell_67_97 ( BL97, BLN97, WL67);
sram_cell_6t_3 inst_cell_67_96 ( BL96, BLN96, WL67);
sram_cell_6t_3 inst_cell_67_95 ( BL95, BLN95, WL67);
sram_cell_6t_3 inst_cell_67_94 ( BL94, BLN94, WL67);
sram_cell_6t_3 inst_cell_67_93 ( BL93, BLN93, WL67);
sram_cell_6t_3 inst_cell_67_92 ( BL92, BLN92, WL67);
sram_cell_6t_3 inst_cell_67_91 ( BL91, BLN91, WL67);
sram_cell_6t_3 inst_cell_67_90 ( BL90, BLN90, WL67);
sram_cell_6t_3 inst_cell_67_89 ( BL89, BLN89, WL67);
sram_cell_6t_3 inst_cell_67_88 ( BL88, BLN88, WL67);
sram_cell_6t_3 inst_cell_67_87 ( BL87, BLN87, WL67);
sram_cell_6t_3 inst_cell_67_86 ( BL86, BLN86, WL67);
sram_cell_6t_3 inst_cell_67_85 ( BL85, BLN85, WL67);
sram_cell_6t_3 inst_cell_67_84 ( BL84, BLN84, WL67);
sram_cell_6t_3 inst_cell_67_83 ( BL83, BLN83, WL67);
sram_cell_6t_3 inst_cell_67_82 ( BL82, BLN82, WL67);
sram_cell_6t_3 inst_cell_67_81 ( BL81, BLN81, WL67);
sram_cell_6t_3 inst_cell_67_80 ( BL80, BLN80, WL67);
sram_cell_6t_3 inst_cell_67_79 ( BL79, BLN79, WL67);
sram_cell_6t_3 inst_cell_67_78 ( BL78, BLN78, WL67);
sram_cell_6t_3 inst_cell_67_77 ( BL77, BLN77, WL67);
sram_cell_6t_3 inst_cell_67_76 ( BL76, BLN76, WL67);
sram_cell_6t_3 inst_cell_67_75 ( BL75, BLN75, WL67);
sram_cell_6t_3 inst_cell_67_74 ( BL74, BLN74, WL67);
sram_cell_6t_3 inst_cell_67_73 ( BL73, BLN73, WL67);
sram_cell_6t_3 inst_cell_67_72 ( BL72, BLN72, WL67);
sram_cell_6t_3 inst_cell_67_71 ( BL71, BLN71, WL67);
sram_cell_6t_3 inst_cell_67_70 ( BL70, BLN70, WL67);
sram_cell_6t_3 inst_cell_67_69 ( BL69, BLN69, WL67);
sram_cell_6t_3 inst_cell_67_68 ( BL68, BLN68, WL67);
sram_cell_6t_3 inst_cell_67_67 ( BL67, BLN67, WL67);
sram_cell_6t_3 inst_cell_67_66 ( BL66, BLN66, WL67);
sram_cell_6t_3 inst_cell_67_65 ( BL65, BLN65, WL67);
sram_cell_6t_3 inst_cell_67_64 ( BL64, BLN64, WL67);
sram_cell_6t_3 inst_cell_67_63 ( BL63, BLN63, WL67);
sram_cell_6t_3 inst_cell_67_62 ( BL62, BLN62, WL67);
sram_cell_6t_3 inst_cell_67_61 ( BL61, BLN61, WL67);
sram_cell_6t_3 inst_cell_67_60 ( BL60, BLN60, WL67);
sram_cell_6t_3 inst_cell_67_59 ( BL59, BLN59, WL67);
sram_cell_6t_3 inst_cell_67_58 ( BL58, BLN58, WL67);
sram_cell_6t_3 inst_cell_67_57 ( BL57, BLN57, WL67);
sram_cell_6t_3 inst_cell_67_56 ( BL56, BLN56, WL67);
sram_cell_6t_3 inst_cell_67_55 ( BL55, BLN55, WL67);
sram_cell_6t_3 inst_cell_67_54 ( BL54, BLN54, WL67);
sram_cell_6t_3 inst_cell_67_53 ( BL53, BLN53, WL67);
sram_cell_6t_3 inst_cell_67_52 ( BL52, BLN52, WL67);
sram_cell_6t_3 inst_cell_67_51 ( BL51, BLN51, WL67);
sram_cell_6t_3 inst_cell_67_50 ( BL50, BLN50, WL67);
sram_cell_6t_3 inst_cell_67_49 ( BL49, BLN49, WL67);
sram_cell_6t_3 inst_cell_67_48 ( BL48, BLN48, WL67);
sram_cell_6t_3 inst_cell_67_47 ( BL47, BLN47, WL67);
sram_cell_6t_3 inst_cell_67_46 ( BL46, BLN46, WL67);
sram_cell_6t_3 inst_cell_67_45 ( BL45, BLN45, WL67);
sram_cell_6t_3 inst_cell_67_44 ( BL44, BLN44, WL67);
sram_cell_6t_3 inst_cell_67_43 ( BL43, BLN43, WL67);
sram_cell_6t_3 inst_cell_67_42 ( BL42, BLN42, WL67);
sram_cell_6t_3 inst_cell_67_41 ( BL41, BLN41, WL67);
sram_cell_6t_3 inst_cell_67_40 ( BL40, BLN40, WL67);
sram_cell_6t_3 inst_cell_67_39 ( BL39, BLN39, WL67);
sram_cell_6t_3 inst_cell_67_38 ( BL38, BLN38, WL67);
sram_cell_6t_3 inst_cell_67_37 ( BL37, BLN37, WL67);
sram_cell_6t_3 inst_cell_67_36 ( BL36, BLN36, WL67);
sram_cell_6t_3 inst_cell_67_35 ( BL35, BLN35, WL67);
sram_cell_6t_3 inst_cell_67_34 ( BL34, BLN34, WL67);
sram_cell_6t_3 inst_cell_67_33 ( BL33, BLN33, WL67);
sram_cell_6t_3 inst_cell_67_32 ( BL32, BLN32, WL67);
sram_cell_6t_3 inst_cell_67_31 ( BL31, BLN31, WL67);
sram_cell_6t_3 inst_cell_67_30 ( BL30, BLN30, WL67);
sram_cell_6t_3 inst_cell_67_29 ( BL29, BLN29, WL67);
sram_cell_6t_3 inst_cell_67_28 ( BL28, BLN28, WL67);
sram_cell_6t_3 inst_cell_67_27 ( BL27, BLN27, WL67);
sram_cell_6t_3 inst_cell_67_26 ( BL26, BLN26, WL67);
sram_cell_6t_3 inst_cell_67_25 ( BL25, BLN25, WL67);
sram_cell_6t_3 inst_cell_67_24 ( BL24, BLN24, WL67);
sram_cell_6t_3 inst_cell_67_23 ( BL23, BLN23, WL67);
sram_cell_6t_3 inst_cell_67_22 ( BL22, BLN22, WL67);
sram_cell_6t_3 inst_cell_67_21 ( BL21, BLN21, WL67);
sram_cell_6t_3 inst_cell_67_20 ( BL20, BLN20, WL67);
sram_cell_6t_3 inst_cell_67_19 ( BL19, BLN19, WL67);
sram_cell_6t_3 inst_cell_67_18 ( BL18, BLN18, WL67);
sram_cell_6t_3 inst_cell_67_17 ( BL17, BLN17, WL67);
sram_cell_6t_3 inst_cell_67_16 ( BL16, BLN16, WL67);
sram_cell_6t_3 inst_cell_67_15 ( BL15, BLN15, WL67);
sram_cell_6t_3 inst_cell_67_14 ( BL14, BLN14, WL67);
sram_cell_6t_3 inst_cell_67_13 ( BL13, BLN13, WL67);
sram_cell_6t_3 inst_cell_67_12 ( BL12, BLN12, WL67);
sram_cell_6t_3 inst_cell_67_11 ( BL11, BLN11, WL67);
sram_cell_6t_3 inst_cell_67_10 ( BL10, BLN10, WL67);
sram_cell_6t_3 inst_cell_67_9 ( BL9, BLN9, WL67);
sram_cell_6t_3 inst_cell_67_8 ( BL8, BLN8, WL67);
sram_cell_6t_3 inst_cell_67_7 ( BL7, BLN7, WL67);
sram_cell_6t_3 inst_cell_67_6 ( BL6, BLN6, WL67);
sram_cell_6t_3 inst_cell_67_5 ( BL5, BLN5, WL67);
sram_cell_6t_3 inst_cell_67_4 ( BL4, BLN4, WL67);
sram_cell_6t_3 inst_cell_67_3 ( BL3, BLN3, WL67);
sram_cell_6t_3 inst_cell_67_2 ( BL2, BLN2, WL67);
sram_cell_6t_3 inst_cell_67_1 ( BL1, BLN1, WL67);
sram_cell_6t_3 inst_cell_67_0 ( BL0, BLN0, WL67);
sram_cell_6t_3 inst_cell_66_127 ( BL127, BLN127, WL66);
sram_cell_6t_3 inst_cell_66_126 ( BL126, BLN126, WL66);
sram_cell_6t_3 inst_cell_66_125 ( BL125, BLN125, WL66);
sram_cell_6t_3 inst_cell_66_124 ( BL124, BLN124, WL66);
sram_cell_6t_3 inst_cell_66_123 ( BL123, BLN123, WL66);
sram_cell_6t_3 inst_cell_66_122 ( BL122, BLN122, WL66);
sram_cell_6t_3 inst_cell_66_121 ( BL121, BLN121, WL66);
sram_cell_6t_3 inst_cell_66_120 ( BL120, BLN120, WL66);
sram_cell_6t_3 inst_cell_66_119 ( BL119, BLN119, WL66);
sram_cell_6t_3 inst_cell_66_118 ( BL118, BLN118, WL66);
sram_cell_6t_3 inst_cell_66_117 ( BL117, BLN117, WL66);
sram_cell_6t_3 inst_cell_66_116 ( BL116, BLN116, WL66);
sram_cell_6t_3 inst_cell_66_115 ( BL115, BLN115, WL66);
sram_cell_6t_3 inst_cell_66_114 ( BL114, BLN114, WL66);
sram_cell_6t_3 inst_cell_66_113 ( BL113, BLN113, WL66);
sram_cell_6t_3 inst_cell_66_112 ( BL112, BLN112, WL66);
sram_cell_6t_3 inst_cell_66_111 ( BL111, BLN111, WL66);
sram_cell_6t_3 inst_cell_66_110 ( BL110, BLN110, WL66);
sram_cell_6t_3 inst_cell_66_109 ( BL109, BLN109, WL66);
sram_cell_6t_3 inst_cell_66_108 ( BL108, BLN108, WL66);
sram_cell_6t_3 inst_cell_66_107 ( BL107, BLN107, WL66);
sram_cell_6t_3 inst_cell_66_106 ( BL106, BLN106, WL66);
sram_cell_6t_3 inst_cell_66_105 ( BL105, BLN105, WL66);
sram_cell_6t_3 inst_cell_66_104 ( BL104, BLN104, WL66);
sram_cell_6t_3 inst_cell_66_103 ( BL103, BLN103, WL66);
sram_cell_6t_3 inst_cell_66_102 ( BL102, BLN102, WL66);
sram_cell_6t_3 inst_cell_66_101 ( BL101, BLN101, WL66);
sram_cell_6t_3 inst_cell_66_100 ( BL100, BLN100, WL66);
sram_cell_6t_3 inst_cell_66_99 ( BL99, BLN99, WL66);
sram_cell_6t_3 inst_cell_66_98 ( BL98, BLN98, WL66);
sram_cell_6t_3 inst_cell_66_97 ( BL97, BLN97, WL66);
sram_cell_6t_3 inst_cell_66_96 ( BL96, BLN96, WL66);
sram_cell_6t_3 inst_cell_66_95 ( BL95, BLN95, WL66);
sram_cell_6t_3 inst_cell_66_94 ( BL94, BLN94, WL66);
sram_cell_6t_3 inst_cell_66_93 ( BL93, BLN93, WL66);
sram_cell_6t_3 inst_cell_66_92 ( BL92, BLN92, WL66);
sram_cell_6t_3 inst_cell_66_91 ( BL91, BLN91, WL66);
sram_cell_6t_3 inst_cell_66_90 ( BL90, BLN90, WL66);
sram_cell_6t_3 inst_cell_66_89 ( BL89, BLN89, WL66);
sram_cell_6t_3 inst_cell_66_88 ( BL88, BLN88, WL66);
sram_cell_6t_3 inst_cell_66_87 ( BL87, BLN87, WL66);
sram_cell_6t_3 inst_cell_66_86 ( BL86, BLN86, WL66);
sram_cell_6t_3 inst_cell_66_85 ( BL85, BLN85, WL66);
sram_cell_6t_3 inst_cell_66_84 ( BL84, BLN84, WL66);
sram_cell_6t_3 inst_cell_66_83 ( BL83, BLN83, WL66);
sram_cell_6t_3 inst_cell_66_82 ( BL82, BLN82, WL66);
sram_cell_6t_3 inst_cell_66_81 ( BL81, BLN81, WL66);
sram_cell_6t_3 inst_cell_66_80 ( BL80, BLN80, WL66);
sram_cell_6t_3 inst_cell_66_79 ( BL79, BLN79, WL66);
sram_cell_6t_3 inst_cell_66_78 ( BL78, BLN78, WL66);
sram_cell_6t_3 inst_cell_66_77 ( BL77, BLN77, WL66);
sram_cell_6t_3 inst_cell_66_76 ( BL76, BLN76, WL66);
sram_cell_6t_3 inst_cell_66_75 ( BL75, BLN75, WL66);
sram_cell_6t_3 inst_cell_66_74 ( BL74, BLN74, WL66);
sram_cell_6t_3 inst_cell_66_73 ( BL73, BLN73, WL66);
sram_cell_6t_3 inst_cell_66_72 ( BL72, BLN72, WL66);
sram_cell_6t_3 inst_cell_66_71 ( BL71, BLN71, WL66);
sram_cell_6t_3 inst_cell_66_70 ( BL70, BLN70, WL66);
sram_cell_6t_3 inst_cell_66_69 ( BL69, BLN69, WL66);
sram_cell_6t_3 inst_cell_66_68 ( BL68, BLN68, WL66);
sram_cell_6t_3 inst_cell_66_67 ( BL67, BLN67, WL66);
sram_cell_6t_3 inst_cell_66_66 ( BL66, BLN66, WL66);
sram_cell_6t_3 inst_cell_66_65 ( BL65, BLN65, WL66);
sram_cell_6t_3 inst_cell_66_64 ( BL64, BLN64, WL66);
sram_cell_6t_3 inst_cell_66_63 ( BL63, BLN63, WL66);
sram_cell_6t_3 inst_cell_66_62 ( BL62, BLN62, WL66);
sram_cell_6t_3 inst_cell_66_61 ( BL61, BLN61, WL66);
sram_cell_6t_3 inst_cell_66_60 ( BL60, BLN60, WL66);
sram_cell_6t_3 inst_cell_66_59 ( BL59, BLN59, WL66);
sram_cell_6t_3 inst_cell_66_58 ( BL58, BLN58, WL66);
sram_cell_6t_3 inst_cell_66_57 ( BL57, BLN57, WL66);
sram_cell_6t_3 inst_cell_66_56 ( BL56, BLN56, WL66);
sram_cell_6t_3 inst_cell_66_55 ( BL55, BLN55, WL66);
sram_cell_6t_3 inst_cell_66_54 ( BL54, BLN54, WL66);
sram_cell_6t_3 inst_cell_66_53 ( BL53, BLN53, WL66);
sram_cell_6t_3 inst_cell_66_52 ( BL52, BLN52, WL66);
sram_cell_6t_3 inst_cell_66_51 ( BL51, BLN51, WL66);
sram_cell_6t_3 inst_cell_66_50 ( BL50, BLN50, WL66);
sram_cell_6t_3 inst_cell_66_49 ( BL49, BLN49, WL66);
sram_cell_6t_3 inst_cell_66_48 ( BL48, BLN48, WL66);
sram_cell_6t_3 inst_cell_66_47 ( BL47, BLN47, WL66);
sram_cell_6t_3 inst_cell_66_46 ( BL46, BLN46, WL66);
sram_cell_6t_3 inst_cell_66_45 ( BL45, BLN45, WL66);
sram_cell_6t_3 inst_cell_66_44 ( BL44, BLN44, WL66);
sram_cell_6t_3 inst_cell_66_43 ( BL43, BLN43, WL66);
sram_cell_6t_3 inst_cell_66_42 ( BL42, BLN42, WL66);
sram_cell_6t_3 inst_cell_66_41 ( BL41, BLN41, WL66);
sram_cell_6t_3 inst_cell_66_40 ( BL40, BLN40, WL66);
sram_cell_6t_3 inst_cell_66_39 ( BL39, BLN39, WL66);
sram_cell_6t_3 inst_cell_66_38 ( BL38, BLN38, WL66);
sram_cell_6t_3 inst_cell_66_37 ( BL37, BLN37, WL66);
sram_cell_6t_3 inst_cell_66_36 ( BL36, BLN36, WL66);
sram_cell_6t_3 inst_cell_66_35 ( BL35, BLN35, WL66);
sram_cell_6t_3 inst_cell_66_34 ( BL34, BLN34, WL66);
sram_cell_6t_3 inst_cell_66_33 ( BL33, BLN33, WL66);
sram_cell_6t_3 inst_cell_66_32 ( BL32, BLN32, WL66);
sram_cell_6t_3 inst_cell_66_31 ( BL31, BLN31, WL66);
sram_cell_6t_3 inst_cell_66_30 ( BL30, BLN30, WL66);
sram_cell_6t_3 inst_cell_66_29 ( BL29, BLN29, WL66);
sram_cell_6t_3 inst_cell_66_28 ( BL28, BLN28, WL66);
sram_cell_6t_3 inst_cell_66_27 ( BL27, BLN27, WL66);
sram_cell_6t_3 inst_cell_66_26 ( BL26, BLN26, WL66);
sram_cell_6t_3 inst_cell_66_25 ( BL25, BLN25, WL66);
sram_cell_6t_3 inst_cell_66_24 ( BL24, BLN24, WL66);
sram_cell_6t_3 inst_cell_66_23 ( BL23, BLN23, WL66);
sram_cell_6t_3 inst_cell_66_22 ( BL22, BLN22, WL66);
sram_cell_6t_3 inst_cell_66_21 ( BL21, BLN21, WL66);
sram_cell_6t_3 inst_cell_66_20 ( BL20, BLN20, WL66);
sram_cell_6t_3 inst_cell_66_19 ( BL19, BLN19, WL66);
sram_cell_6t_3 inst_cell_66_18 ( BL18, BLN18, WL66);
sram_cell_6t_3 inst_cell_66_17 ( BL17, BLN17, WL66);
sram_cell_6t_3 inst_cell_66_16 ( BL16, BLN16, WL66);
sram_cell_6t_3 inst_cell_66_15 ( BL15, BLN15, WL66);
sram_cell_6t_3 inst_cell_66_14 ( BL14, BLN14, WL66);
sram_cell_6t_3 inst_cell_66_13 ( BL13, BLN13, WL66);
sram_cell_6t_3 inst_cell_66_12 ( BL12, BLN12, WL66);
sram_cell_6t_3 inst_cell_66_11 ( BL11, BLN11, WL66);
sram_cell_6t_3 inst_cell_66_10 ( BL10, BLN10, WL66);
sram_cell_6t_3 inst_cell_66_9 ( BL9, BLN9, WL66);
sram_cell_6t_3 inst_cell_66_8 ( BL8, BLN8, WL66);
sram_cell_6t_3 inst_cell_66_7 ( BL7, BLN7, WL66);
sram_cell_6t_3 inst_cell_66_6 ( BL6, BLN6, WL66);
sram_cell_6t_3 inst_cell_66_5 ( BL5, BLN5, WL66);
sram_cell_6t_3 inst_cell_66_4 ( BL4, BLN4, WL66);
sram_cell_6t_3 inst_cell_66_3 ( BL3, BLN3, WL66);
sram_cell_6t_3 inst_cell_66_2 ( BL2, BLN2, WL66);
sram_cell_6t_3 inst_cell_66_1 ( BL1, BLN1, WL66);
sram_cell_6t_3 inst_cell_66_0 ( BL0, BLN0, WL66);
sram_cell_6t_3 inst_cell_65_127 ( BL127, BLN127, WL65);
sram_cell_6t_3 inst_cell_65_126 ( BL126, BLN126, WL65);
sram_cell_6t_3 inst_cell_65_125 ( BL125, BLN125, WL65);
sram_cell_6t_3 inst_cell_65_124 ( BL124, BLN124, WL65);
sram_cell_6t_3 inst_cell_65_123 ( BL123, BLN123, WL65);
sram_cell_6t_3 inst_cell_65_122 ( BL122, BLN122, WL65);
sram_cell_6t_3 inst_cell_65_121 ( BL121, BLN121, WL65);
sram_cell_6t_3 inst_cell_65_120 ( BL120, BLN120, WL65);
sram_cell_6t_3 inst_cell_65_119 ( BL119, BLN119, WL65);
sram_cell_6t_3 inst_cell_65_118 ( BL118, BLN118, WL65);
sram_cell_6t_3 inst_cell_65_117 ( BL117, BLN117, WL65);
sram_cell_6t_3 inst_cell_65_116 ( BL116, BLN116, WL65);
sram_cell_6t_3 inst_cell_65_115 ( BL115, BLN115, WL65);
sram_cell_6t_3 inst_cell_65_114 ( BL114, BLN114, WL65);
sram_cell_6t_3 inst_cell_65_113 ( BL113, BLN113, WL65);
sram_cell_6t_3 inst_cell_65_112 ( BL112, BLN112, WL65);
sram_cell_6t_3 inst_cell_65_111 ( BL111, BLN111, WL65);
sram_cell_6t_3 inst_cell_65_110 ( BL110, BLN110, WL65);
sram_cell_6t_3 inst_cell_65_109 ( BL109, BLN109, WL65);
sram_cell_6t_3 inst_cell_65_108 ( BL108, BLN108, WL65);
sram_cell_6t_3 inst_cell_65_107 ( BL107, BLN107, WL65);
sram_cell_6t_3 inst_cell_65_106 ( BL106, BLN106, WL65);
sram_cell_6t_3 inst_cell_65_105 ( BL105, BLN105, WL65);
sram_cell_6t_3 inst_cell_65_104 ( BL104, BLN104, WL65);
sram_cell_6t_3 inst_cell_65_103 ( BL103, BLN103, WL65);
sram_cell_6t_3 inst_cell_65_102 ( BL102, BLN102, WL65);
sram_cell_6t_3 inst_cell_65_101 ( BL101, BLN101, WL65);
sram_cell_6t_3 inst_cell_65_100 ( BL100, BLN100, WL65);
sram_cell_6t_3 inst_cell_65_99 ( BL99, BLN99, WL65);
sram_cell_6t_3 inst_cell_65_98 ( BL98, BLN98, WL65);
sram_cell_6t_3 inst_cell_65_97 ( BL97, BLN97, WL65);
sram_cell_6t_3 inst_cell_65_96 ( BL96, BLN96, WL65);
sram_cell_6t_3 inst_cell_65_95 ( BL95, BLN95, WL65);
sram_cell_6t_3 inst_cell_65_94 ( BL94, BLN94, WL65);
sram_cell_6t_3 inst_cell_65_93 ( BL93, BLN93, WL65);
sram_cell_6t_3 inst_cell_65_92 ( BL92, BLN92, WL65);
sram_cell_6t_3 inst_cell_65_91 ( BL91, BLN91, WL65);
sram_cell_6t_3 inst_cell_65_90 ( BL90, BLN90, WL65);
sram_cell_6t_3 inst_cell_65_89 ( BL89, BLN89, WL65);
sram_cell_6t_3 inst_cell_65_88 ( BL88, BLN88, WL65);
sram_cell_6t_3 inst_cell_65_87 ( BL87, BLN87, WL65);
sram_cell_6t_3 inst_cell_65_86 ( BL86, BLN86, WL65);
sram_cell_6t_3 inst_cell_65_85 ( BL85, BLN85, WL65);
sram_cell_6t_3 inst_cell_65_84 ( BL84, BLN84, WL65);
sram_cell_6t_3 inst_cell_65_83 ( BL83, BLN83, WL65);
sram_cell_6t_3 inst_cell_65_82 ( BL82, BLN82, WL65);
sram_cell_6t_3 inst_cell_65_81 ( BL81, BLN81, WL65);
sram_cell_6t_3 inst_cell_65_80 ( BL80, BLN80, WL65);
sram_cell_6t_3 inst_cell_65_79 ( BL79, BLN79, WL65);
sram_cell_6t_3 inst_cell_65_78 ( BL78, BLN78, WL65);
sram_cell_6t_3 inst_cell_65_77 ( BL77, BLN77, WL65);
sram_cell_6t_3 inst_cell_65_76 ( BL76, BLN76, WL65);
sram_cell_6t_3 inst_cell_65_75 ( BL75, BLN75, WL65);
sram_cell_6t_3 inst_cell_65_74 ( BL74, BLN74, WL65);
sram_cell_6t_3 inst_cell_65_73 ( BL73, BLN73, WL65);
sram_cell_6t_3 inst_cell_65_72 ( BL72, BLN72, WL65);
sram_cell_6t_3 inst_cell_65_71 ( BL71, BLN71, WL65);
sram_cell_6t_3 inst_cell_65_70 ( BL70, BLN70, WL65);
sram_cell_6t_3 inst_cell_65_69 ( BL69, BLN69, WL65);
sram_cell_6t_3 inst_cell_65_68 ( BL68, BLN68, WL65);
sram_cell_6t_3 inst_cell_65_67 ( BL67, BLN67, WL65);
sram_cell_6t_3 inst_cell_65_66 ( BL66, BLN66, WL65);
sram_cell_6t_3 inst_cell_65_65 ( BL65, BLN65, WL65);
sram_cell_6t_3 inst_cell_65_64 ( BL64, BLN64, WL65);
sram_cell_6t_3 inst_cell_65_63 ( BL63, BLN63, WL65);
sram_cell_6t_3 inst_cell_65_62 ( BL62, BLN62, WL65);
sram_cell_6t_3 inst_cell_65_61 ( BL61, BLN61, WL65);
sram_cell_6t_3 inst_cell_65_60 ( BL60, BLN60, WL65);
sram_cell_6t_3 inst_cell_65_59 ( BL59, BLN59, WL65);
sram_cell_6t_3 inst_cell_65_58 ( BL58, BLN58, WL65);
sram_cell_6t_3 inst_cell_65_57 ( BL57, BLN57, WL65);
sram_cell_6t_3 inst_cell_65_56 ( BL56, BLN56, WL65);
sram_cell_6t_3 inst_cell_65_55 ( BL55, BLN55, WL65);
sram_cell_6t_3 inst_cell_65_54 ( BL54, BLN54, WL65);
sram_cell_6t_3 inst_cell_65_53 ( BL53, BLN53, WL65);
sram_cell_6t_3 inst_cell_65_52 ( BL52, BLN52, WL65);
sram_cell_6t_3 inst_cell_65_51 ( BL51, BLN51, WL65);
sram_cell_6t_3 inst_cell_65_50 ( BL50, BLN50, WL65);
sram_cell_6t_3 inst_cell_65_49 ( BL49, BLN49, WL65);
sram_cell_6t_3 inst_cell_65_48 ( BL48, BLN48, WL65);
sram_cell_6t_3 inst_cell_65_47 ( BL47, BLN47, WL65);
sram_cell_6t_3 inst_cell_65_46 ( BL46, BLN46, WL65);
sram_cell_6t_3 inst_cell_65_45 ( BL45, BLN45, WL65);
sram_cell_6t_3 inst_cell_65_44 ( BL44, BLN44, WL65);
sram_cell_6t_3 inst_cell_65_43 ( BL43, BLN43, WL65);
sram_cell_6t_3 inst_cell_65_42 ( BL42, BLN42, WL65);
sram_cell_6t_3 inst_cell_65_41 ( BL41, BLN41, WL65);
sram_cell_6t_3 inst_cell_65_40 ( BL40, BLN40, WL65);
sram_cell_6t_3 inst_cell_65_39 ( BL39, BLN39, WL65);
sram_cell_6t_3 inst_cell_65_38 ( BL38, BLN38, WL65);
sram_cell_6t_3 inst_cell_65_37 ( BL37, BLN37, WL65);
sram_cell_6t_3 inst_cell_65_36 ( BL36, BLN36, WL65);
sram_cell_6t_3 inst_cell_65_35 ( BL35, BLN35, WL65);
sram_cell_6t_3 inst_cell_65_34 ( BL34, BLN34, WL65);
sram_cell_6t_3 inst_cell_65_33 ( BL33, BLN33, WL65);
sram_cell_6t_3 inst_cell_65_32 ( BL32, BLN32, WL65);
sram_cell_6t_3 inst_cell_65_31 ( BL31, BLN31, WL65);
sram_cell_6t_3 inst_cell_65_30 ( BL30, BLN30, WL65);
sram_cell_6t_3 inst_cell_65_29 ( BL29, BLN29, WL65);
sram_cell_6t_3 inst_cell_65_28 ( BL28, BLN28, WL65);
sram_cell_6t_3 inst_cell_65_27 ( BL27, BLN27, WL65);
sram_cell_6t_3 inst_cell_65_26 ( BL26, BLN26, WL65);
sram_cell_6t_3 inst_cell_65_25 ( BL25, BLN25, WL65);
sram_cell_6t_3 inst_cell_65_24 ( BL24, BLN24, WL65);
sram_cell_6t_3 inst_cell_65_23 ( BL23, BLN23, WL65);
sram_cell_6t_3 inst_cell_65_22 ( BL22, BLN22, WL65);
sram_cell_6t_3 inst_cell_65_21 ( BL21, BLN21, WL65);
sram_cell_6t_3 inst_cell_65_20 ( BL20, BLN20, WL65);
sram_cell_6t_3 inst_cell_65_19 ( BL19, BLN19, WL65);
sram_cell_6t_3 inst_cell_65_18 ( BL18, BLN18, WL65);
sram_cell_6t_3 inst_cell_65_17 ( BL17, BLN17, WL65);
sram_cell_6t_3 inst_cell_65_16 ( BL16, BLN16, WL65);
sram_cell_6t_3 inst_cell_65_15 ( BL15, BLN15, WL65);
sram_cell_6t_3 inst_cell_65_14 ( BL14, BLN14, WL65);
sram_cell_6t_3 inst_cell_65_13 ( BL13, BLN13, WL65);
sram_cell_6t_3 inst_cell_65_12 ( BL12, BLN12, WL65);
sram_cell_6t_3 inst_cell_65_11 ( BL11, BLN11, WL65);
sram_cell_6t_3 inst_cell_65_10 ( BL10, BLN10, WL65);
sram_cell_6t_3 inst_cell_65_9 ( BL9, BLN9, WL65);
sram_cell_6t_3 inst_cell_65_8 ( BL8, BLN8, WL65);
sram_cell_6t_3 inst_cell_65_7 ( BL7, BLN7, WL65);
sram_cell_6t_3 inst_cell_65_6 ( BL6, BLN6, WL65);
sram_cell_6t_3 inst_cell_65_5 ( BL5, BLN5, WL65);
sram_cell_6t_3 inst_cell_65_4 ( BL4, BLN4, WL65);
sram_cell_6t_3 inst_cell_65_3 ( BL3, BLN3, WL65);
sram_cell_6t_3 inst_cell_65_2 ( BL2, BLN2, WL65);
sram_cell_6t_3 inst_cell_65_1 ( BL1, BLN1, WL65);
sram_cell_6t_3 inst_cell_65_0 ( BL0, BLN0, WL65);
sram_cell_6t_3 inst_cell_64_127 ( BL127, BLN127, WL64);
sram_cell_6t_3 inst_cell_64_126 ( BL126, BLN126, WL64);
sram_cell_6t_3 inst_cell_64_125 ( BL125, BLN125, WL64);
sram_cell_6t_3 inst_cell_64_124 ( BL124, BLN124, WL64);
sram_cell_6t_3 inst_cell_64_123 ( BL123, BLN123, WL64);
sram_cell_6t_3 inst_cell_64_122 ( BL122, BLN122, WL64);
sram_cell_6t_3 inst_cell_64_121 ( BL121, BLN121, WL64);
sram_cell_6t_3 inst_cell_64_120 ( BL120, BLN120, WL64);
sram_cell_6t_3 inst_cell_64_119 ( BL119, BLN119, WL64);
sram_cell_6t_3 inst_cell_64_118 ( BL118, BLN118, WL64);
sram_cell_6t_3 inst_cell_64_117 ( BL117, BLN117, WL64);
sram_cell_6t_3 inst_cell_64_116 ( BL116, BLN116, WL64);
sram_cell_6t_3 inst_cell_64_115 ( BL115, BLN115, WL64);
sram_cell_6t_3 inst_cell_64_114 ( BL114, BLN114, WL64);
sram_cell_6t_3 inst_cell_64_113 ( BL113, BLN113, WL64);
sram_cell_6t_3 inst_cell_64_112 ( BL112, BLN112, WL64);
sram_cell_6t_3 inst_cell_64_111 ( BL111, BLN111, WL64);
sram_cell_6t_3 inst_cell_64_110 ( BL110, BLN110, WL64);
sram_cell_6t_3 inst_cell_64_109 ( BL109, BLN109, WL64);
sram_cell_6t_3 inst_cell_64_108 ( BL108, BLN108, WL64);
sram_cell_6t_3 inst_cell_64_107 ( BL107, BLN107, WL64);
sram_cell_6t_3 inst_cell_64_106 ( BL106, BLN106, WL64);
sram_cell_6t_3 inst_cell_64_105 ( BL105, BLN105, WL64);
sram_cell_6t_3 inst_cell_64_104 ( BL104, BLN104, WL64);
sram_cell_6t_3 inst_cell_64_103 ( BL103, BLN103, WL64);
sram_cell_6t_3 inst_cell_64_102 ( BL102, BLN102, WL64);
sram_cell_6t_3 inst_cell_64_101 ( BL101, BLN101, WL64);
sram_cell_6t_3 inst_cell_64_100 ( BL100, BLN100, WL64);
sram_cell_6t_3 inst_cell_64_99 ( BL99, BLN99, WL64);
sram_cell_6t_3 inst_cell_64_98 ( BL98, BLN98, WL64);
sram_cell_6t_3 inst_cell_64_97 ( BL97, BLN97, WL64);
sram_cell_6t_3 inst_cell_64_96 ( BL96, BLN96, WL64);
sram_cell_6t_3 inst_cell_64_95 ( BL95, BLN95, WL64);
sram_cell_6t_3 inst_cell_64_94 ( BL94, BLN94, WL64);
sram_cell_6t_3 inst_cell_64_93 ( BL93, BLN93, WL64);
sram_cell_6t_3 inst_cell_64_92 ( BL92, BLN92, WL64);
sram_cell_6t_3 inst_cell_64_91 ( BL91, BLN91, WL64);
sram_cell_6t_3 inst_cell_64_90 ( BL90, BLN90, WL64);
sram_cell_6t_3 inst_cell_64_89 ( BL89, BLN89, WL64);
sram_cell_6t_3 inst_cell_64_88 ( BL88, BLN88, WL64);
sram_cell_6t_3 inst_cell_64_87 ( BL87, BLN87, WL64);
sram_cell_6t_3 inst_cell_64_86 ( BL86, BLN86, WL64);
sram_cell_6t_3 inst_cell_64_85 ( BL85, BLN85, WL64);
sram_cell_6t_3 inst_cell_64_84 ( BL84, BLN84, WL64);
sram_cell_6t_3 inst_cell_64_83 ( BL83, BLN83, WL64);
sram_cell_6t_3 inst_cell_64_82 ( BL82, BLN82, WL64);
sram_cell_6t_3 inst_cell_64_81 ( BL81, BLN81, WL64);
sram_cell_6t_3 inst_cell_64_80 ( BL80, BLN80, WL64);
sram_cell_6t_3 inst_cell_64_79 ( BL79, BLN79, WL64);
sram_cell_6t_3 inst_cell_64_78 ( BL78, BLN78, WL64);
sram_cell_6t_3 inst_cell_64_77 ( BL77, BLN77, WL64);
sram_cell_6t_3 inst_cell_64_76 ( BL76, BLN76, WL64);
sram_cell_6t_3 inst_cell_64_75 ( BL75, BLN75, WL64);
sram_cell_6t_3 inst_cell_64_74 ( BL74, BLN74, WL64);
sram_cell_6t_3 inst_cell_64_73 ( BL73, BLN73, WL64);
sram_cell_6t_3 inst_cell_64_72 ( BL72, BLN72, WL64);
sram_cell_6t_3 inst_cell_64_71 ( BL71, BLN71, WL64);
sram_cell_6t_3 inst_cell_64_70 ( BL70, BLN70, WL64);
sram_cell_6t_3 inst_cell_64_69 ( BL69, BLN69, WL64);
sram_cell_6t_3 inst_cell_64_68 ( BL68, BLN68, WL64);
sram_cell_6t_3 inst_cell_64_67 ( BL67, BLN67, WL64);
sram_cell_6t_3 inst_cell_64_66 ( BL66, BLN66, WL64);
sram_cell_6t_3 inst_cell_64_65 ( BL65, BLN65, WL64);
sram_cell_6t_3 inst_cell_64_64 ( BL64, BLN64, WL64);
sram_cell_6t_3 inst_cell_64_63 ( BL63, BLN63, WL64);
sram_cell_6t_3 inst_cell_64_62 ( BL62, BLN62, WL64);
sram_cell_6t_3 inst_cell_64_61 ( BL61, BLN61, WL64);
sram_cell_6t_3 inst_cell_64_60 ( BL60, BLN60, WL64);
sram_cell_6t_3 inst_cell_64_59 ( BL59, BLN59, WL64);
sram_cell_6t_3 inst_cell_64_58 ( BL58, BLN58, WL64);
sram_cell_6t_3 inst_cell_64_57 ( BL57, BLN57, WL64);
sram_cell_6t_3 inst_cell_64_56 ( BL56, BLN56, WL64);
sram_cell_6t_3 inst_cell_64_55 ( BL55, BLN55, WL64);
sram_cell_6t_3 inst_cell_64_54 ( BL54, BLN54, WL64);
sram_cell_6t_3 inst_cell_64_53 ( BL53, BLN53, WL64);
sram_cell_6t_3 inst_cell_64_52 ( BL52, BLN52, WL64);
sram_cell_6t_3 inst_cell_64_51 ( BL51, BLN51, WL64);
sram_cell_6t_3 inst_cell_64_50 ( BL50, BLN50, WL64);
sram_cell_6t_3 inst_cell_64_49 ( BL49, BLN49, WL64);
sram_cell_6t_3 inst_cell_64_48 ( BL48, BLN48, WL64);
sram_cell_6t_3 inst_cell_64_47 ( BL47, BLN47, WL64);
sram_cell_6t_3 inst_cell_64_46 ( BL46, BLN46, WL64);
sram_cell_6t_3 inst_cell_64_45 ( BL45, BLN45, WL64);
sram_cell_6t_3 inst_cell_64_44 ( BL44, BLN44, WL64);
sram_cell_6t_3 inst_cell_64_43 ( BL43, BLN43, WL64);
sram_cell_6t_3 inst_cell_64_42 ( BL42, BLN42, WL64);
sram_cell_6t_3 inst_cell_64_41 ( BL41, BLN41, WL64);
sram_cell_6t_3 inst_cell_64_40 ( BL40, BLN40, WL64);
sram_cell_6t_3 inst_cell_64_39 ( BL39, BLN39, WL64);
sram_cell_6t_3 inst_cell_64_38 ( BL38, BLN38, WL64);
sram_cell_6t_3 inst_cell_64_37 ( BL37, BLN37, WL64);
sram_cell_6t_3 inst_cell_64_36 ( BL36, BLN36, WL64);
sram_cell_6t_3 inst_cell_64_35 ( BL35, BLN35, WL64);
sram_cell_6t_3 inst_cell_64_34 ( BL34, BLN34, WL64);
sram_cell_6t_3 inst_cell_64_33 ( BL33, BLN33, WL64);
sram_cell_6t_3 inst_cell_64_32 ( BL32, BLN32, WL64);
sram_cell_6t_3 inst_cell_64_31 ( BL31, BLN31, WL64);
sram_cell_6t_3 inst_cell_64_30 ( BL30, BLN30, WL64);
sram_cell_6t_3 inst_cell_64_29 ( BL29, BLN29, WL64);
sram_cell_6t_3 inst_cell_64_28 ( BL28, BLN28, WL64);
sram_cell_6t_3 inst_cell_64_27 ( BL27, BLN27, WL64);
sram_cell_6t_3 inst_cell_64_26 ( BL26, BLN26, WL64);
sram_cell_6t_3 inst_cell_64_25 ( BL25, BLN25, WL64);
sram_cell_6t_3 inst_cell_64_24 ( BL24, BLN24, WL64);
sram_cell_6t_3 inst_cell_64_23 ( BL23, BLN23, WL64);
sram_cell_6t_3 inst_cell_64_22 ( BL22, BLN22, WL64);
sram_cell_6t_3 inst_cell_64_21 ( BL21, BLN21, WL64);
sram_cell_6t_3 inst_cell_64_20 ( BL20, BLN20, WL64);
sram_cell_6t_3 inst_cell_64_19 ( BL19, BLN19, WL64);
sram_cell_6t_3 inst_cell_64_18 ( BL18, BLN18, WL64);
sram_cell_6t_3 inst_cell_64_17 ( BL17, BLN17, WL64);
sram_cell_6t_3 inst_cell_64_16 ( BL16, BLN16, WL64);
sram_cell_6t_3 inst_cell_64_15 ( BL15, BLN15, WL64);
sram_cell_6t_3 inst_cell_64_14 ( BL14, BLN14, WL64);
sram_cell_6t_3 inst_cell_64_13 ( BL13, BLN13, WL64);
sram_cell_6t_3 inst_cell_64_12 ( BL12, BLN12, WL64);
sram_cell_6t_3 inst_cell_64_11 ( BL11, BLN11, WL64);
sram_cell_6t_3 inst_cell_64_10 ( BL10, BLN10, WL64);
sram_cell_6t_3 inst_cell_64_9 ( BL9, BLN9, WL64);
sram_cell_6t_3 inst_cell_64_8 ( BL8, BLN8, WL64);
sram_cell_6t_3 inst_cell_64_7 ( BL7, BLN7, WL64);
sram_cell_6t_3 inst_cell_64_6 ( BL6, BLN6, WL64);
sram_cell_6t_3 inst_cell_64_5 ( BL5, BLN5, WL64);
sram_cell_6t_3 inst_cell_64_4 ( BL4, BLN4, WL64);
sram_cell_6t_3 inst_cell_64_3 ( BL3, BLN3, WL64);
sram_cell_6t_3 inst_cell_64_2 ( BL2, BLN2, WL64);
sram_cell_6t_3 inst_cell_64_1 ( BL1, BLN1, WL64);
sram_cell_6t_3 inst_cell_64_0 ( BL0, BLN0, WL64);
sram_cell_6t_3 inst_cell_63_127 ( BL127, BLN127, WL63);
sram_cell_6t_3 inst_cell_63_126 ( BL126, BLN126, WL63);
sram_cell_6t_3 inst_cell_63_125 ( BL125, BLN125, WL63);
sram_cell_6t_3 inst_cell_63_124 ( BL124, BLN124, WL63);
sram_cell_6t_3 inst_cell_63_123 ( BL123, BLN123, WL63);
sram_cell_6t_3 inst_cell_63_122 ( BL122, BLN122, WL63);
sram_cell_6t_3 inst_cell_63_121 ( BL121, BLN121, WL63);
sram_cell_6t_3 inst_cell_63_120 ( BL120, BLN120, WL63);
sram_cell_6t_3 inst_cell_63_119 ( BL119, BLN119, WL63);
sram_cell_6t_3 inst_cell_63_118 ( BL118, BLN118, WL63);
sram_cell_6t_3 inst_cell_63_117 ( BL117, BLN117, WL63);
sram_cell_6t_3 inst_cell_63_116 ( BL116, BLN116, WL63);
sram_cell_6t_3 inst_cell_63_115 ( BL115, BLN115, WL63);
sram_cell_6t_3 inst_cell_63_114 ( BL114, BLN114, WL63);
sram_cell_6t_3 inst_cell_63_113 ( BL113, BLN113, WL63);
sram_cell_6t_3 inst_cell_63_112 ( BL112, BLN112, WL63);
sram_cell_6t_3 inst_cell_63_111 ( BL111, BLN111, WL63);
sram_cell_6t_3 inst_cell_63_110 ( BL110, BLN110, WL63);
sram_cell_6t_3 inst_cell_63_109 ( BL109, BLN109, WL63);
sram_cell_6t_3 inst_cell_63_108 ( BL108, BLN108, WL63);
sram_cell_6t_3 inst_cell_63_107 ( BL107, BLN107, WL63);
sram_cell_6t_3 inst_cell_63_106 ( BL106, BLN106, WL63);
sram_cell_6t_3 inst_cell_63_105 ( BL105, BLN105, WL63);
sram_cell_6t_3 inst_cell_63_104 ( BL104, BLN104, WL63);
sram_cell_6t_3 inst_cell_63_103 ( BL103, BLN103, WL63);
sram_cell_6t_3 inst_cell_63_102 ( BL102, BLN102, WL63);
sram_cell_6t_3 inst_cell_63_101 ( BL101, BLN101, WL63);
sram_cell_6t_3 inst_cell_63_100 ( BL100, BLN100, WL63);
sram_cell_6t_3 inst_cell_63_99 ( BL99, BLN99, WL63);
sram_cell_6t_3 inst_cell_63_98 ( BL98, BLN98, WL63);
sram_cell_6t_3 inst_cell_63_97 ( BL97, BLN97, WL63);
sram_cell_6t_3 inst_cell_63_96 ( BL96, BLN96, WL63);
sram_cell_6t_3 inst_cell_63_95 ( BL95, BLN95, WL63);
sram_cell_6t_3 inst_cell_63_94 ( BL94, BLN94, WL63);
sram_cell_6t_3 inst_cell_63_93 ( BL93, BLN93, WL63);
sram_cell_6t_3 inst_cell_63_92 ( BL92, BLN92, WL63);
sram_cell_6t_3 inst_cell_63_91 ( BL91, BLN91, WL63);
sram_cell_6t_3 inst_cell_63_90 ( BL90, BLN90, WL63);
sram_cell_6t_3 inst_cell_63_89 ( BL89, BLN89, WL63);
sram_cell_6t_3 inst_cell_63_88 ( BL88, BLN88, WL63);
sram_cell_6t_3 inst_cell_63_87 ( BL87, BLN87, WL63);
sram_cell_6t_3 inst_cell_63_86 ( BL86, BLN86, WL63);
sram_cell_6t_3 inst_cell_63_85 ( BL85, BLN85, WL63);
sram_cell_6t_3 inst_cell_63_84 ( BL84, BLN84, WL63);
sram_cell_6t_3 inst_cell_63_83 ( BL83, BLN83, WL63);
sram_cell_6t_3 inst_cell_63_82 ( BL82, BLN82, WL63);
sram_cell_6t_3 inst_cell_63_81 ( BL81, BLN81, WL63);
sram_cell_6t_3 inst_cell_63_80 ( BL80, BLN80, WL63);
sram_cell_6t_3 inst_cell_63_79 ( BL79, BLN79, WL63);
sram_cell_6t_3 inst_cell_63_78 ( BL78, BLN78, WL63);
sram_cell_6t_3 inst_cell_63_77 ( BL77, BLN77, WL63);
sram_cell_6t_3 inst_cell_63_76 ( BL76, BLN76, WL63);
sram_cell_6t_3 inst_cell_63_75 ( BL75, BLN75, WL63);
sram_cell_6t_3 inst_cell_63_74 ( BL74, BLN74, WL63);
sram_cell_6t_3 inst_cell_63_73 ( BL73, BLN73, WL63);
sram_cell_6t_3 inst_cell_63_72 ( BL72, BLN72, WL63);
sram_cell_6t_3 inst_cell_63_71 ( BL71, BLN71, WL63);
sram_cell_6t_3 inst_cell_63_70 ( BL70, BLN70, WL63);
sram_cell_6t_3 inst_cell_63_69 ( BL69, BLN69, WL63);
sram_cell_6t_3 inst_cell_63_68 ( BL68, BLN68, WL63);
sram_cell_6t_3 inst_cell_63_67 ( BL67, BLN67, WL63);
sram_cell_6t_3 inst_cell_63_66 ( BL66, BLN66, WL63);
sram_cell_6t_3 inst_cell_63_65 ( BL65, BLN65, WL63);
sram_cell_6t_3 inst_cell_63_64 ( BL64, BLN64, WL63);
sram_cell_6t_3 inst_cell_63_63 ( BL63, BLN63, WL63);
sram_cell_6t_3 inst_cell_63_62 ( BL62, BLN62, WL63);
sram_cell_6t_3 inst_cell_63_61 ( BL61, BLN61, WL63);
sram_cell_6t_3 inst_cell_63_60 ( BL60, BLN60, WL63);
sram_cell_6t_3 inst_cell_63_59 ( BL59, BLN59, WL63);
sram_cell_6t_3 inst_cell_63_58 ( BL58, BLN58, WL63);
sram_cell_6t_3 inst_cell_63_57 ( BL57, BLN57, WL63);
sram_cell_6t_3 inst_cell_63_56 ( BL56, BLN56, WL63);
sram_cell_6t_3 inst_cell_63_55 ( BL55, BLN55, WL63);
sram_cell_6t_3 inst_cell_63_54 ( BL54, BLN54, WL63);
sram_cell_6t_3 inst_cell_63_53 ( BL53, BLN53, WL63);
sram_cell_6t_3 inst_cell_63_52 ( BL52, BLN52, WL63);
sram_cell_6t_3 inst_cell_63_51 ( BL51, BLN51, WL63);
sram_cell_6t_3 inst_cell_63_50 ( BL50, BLN50, WL63);
sram_cell_6t_3 inst_cell_63_49 ( BL49, BLN49, WL63);
sram_cell_6t_3 inst_cell_63_48 ( BL48, BLN48, WL63);
sram_cell_6t_3 inst_cell_63_47 ( BL47, BLN47, WL63);
sram_cell_6t_3 inst_cell_63_46 ( BL46, BLN46, WL63);
sram_cell_6t_3 inst_cell_63_45 ( BL45, BLN45, WL63);
sram_cell_6t_3 inst_cell_63_44 ( BL44, BLN44, WL63);
sram_cell_6t_3 inst_cell_63_43 ( BL43, BLN43, WL63);
sram_cell_6t_3 inst_cell_63_42 ( BL42, BLN42, WL63);
sram_cell_6t_3 inst_cell_63_41 ( BL41, BLN41, WL63);
sram_cell_6t_3 inst_cell_63_40 ( BL40, BLN40, WL63);
sram_cell_6t_3 inst_cell_63_39 ( BL39, BLN39, WL63);
sram_cell_6t_3 inst_cell_63_38 ( BL38, BLN38, WL63);
sram_cell_6t_3 inst_cell_63_37 ( BL37, BLN37, WL63);
sram_cell_6t_3 inst_cell_63_36 ( BL36, BLN36, WL63);
sram_cell_6t_3 inst_cell_63_35 ( BL35, BLN35, WL63);
sram_cell_6t_3 inst_cell_63_34 ( BL34, BLN34, WL63);
sram_cell_6t_3 inst_cell_63_33 ( BL33, BLN33, WL63);
sram_cell_6t_3 inst_cell_63_32 ( BL32, BLN32, WL63);
sram_cell_6t_3 inst_cell_63_31 ( BL31, BLN31, WL63);
sram_cell_6t_3 inst_cell_63_30 ( BL30, BLN30, WL63);
sram_cell_6t_3 inst_cell_63_29 ( BL29, BLN29, WL63);
sram_cell_6t_3 inst_cell_63_28 ( BL28, BLN28, WL63);
sram_cell_6t_3 inst_cell_63_27 ( BL27, BLN27, WL63);
sram_cell_6t_3 inst_cell_63_26 ( BL26, BLN26, WL63);
sram_cell_6t_3 inst_cell_63_25 ( BL25, BLN25, WL63);
sram_cell_6t_3 inst_cell_63_24 ( BL24, BLN24, WL63);
sram_cell_6t_3 inst_cell_63_23 ( BL23, BLN23, WL63);
sram_cell_6t_3 inst_cell_63_22 ( BL22, BLN22, WL63);
sram_cell_6t_3 inst_cell_63_21 ( BL21, BLN21, WL63);
sram_cell_6t_3 inst_cell_63_20 ( BL20, BLN20, WL63);
sram_cell_6t_3 inst_cell_63_19 ( BL19, BLN19, WL63);
sram_cell_6t_3 inst_cell_63_18 ( BL18, BLN18, WL63);
sram_cell_6t_3 inst_cell_63_17 ( BL17, BLN17, WL63);
sram_cell_6t_3 inst_cell_63_16 ( BL16, BLN16, WL63);
sram_cell_6t_3 inst_cell_63_15 ( BL15, BLN15, WL63);
sram_cell_6t_3 inst_cell_63_14 ( BL14, BLN14, WL63);
sram_cell_6t_3 inst_cell_63_13 ( BL13, BLN13, WL63);
sram_cell_6t_3 inst_cell_63_12 ( BL12, BLN12, WL63);
sram_cell_6t_3 inst_cell_63_11 ( BL11, BLN11, WL63);
sram_cell_6t_3 inst_cell_63_10 ( BL10, BLN10, WL63);
sram_cell_6t_3 inst_cell_63_9 ( BL9, BLN9, WL63);
sram_cell_6t_3 inst_cell_63_8 ( BL8, BLN8, WL63);
sram_cell_6t_3 inst_cell_63_7 ( BL7, BLN7, WL63);
sram_cell_6t_3 inst_cell_63_6 ( BL6, BLN6, WL63);
sram_cell_6t_3 inst_cell_63_5 ( BL5, BLN5, WL63);
sram_cell_6t_3 inst_cell_63_4 ( BL4, BLN4, WL63);
sram_cell_6t_3 inst_cell_63_3 ( BL3, BLN3, WL63);
sram_cell_6t_3 inst_cell_63_2 ( BL2, BLN2, WL63);
sram_cell_6t_3 inst_cell_63_1 ( BL1, BLN1, WL63);
sram_cell_6t_3 inst_cell_63_0 ( BL0, BLN0, WL63);
sram_cell_6t_3 inst_cell_62_127 ( BL127, BLN127, WL62);
sram_cell_6t_3 inst_cell_62_126 ( BL126, BLN126, WL62);
sram_cell_6t_3 inst_cell_62_125 ( BL125, BLN125, WL62);
sram_cell_6t_3 inst_cell_62_124 ( BL124, BLN124, WL62);
sram_cell_6t_3 inst_cell_62_123 ( BL123, BLN123, WL62);
sram_cell_6t_3 inst_cell_62_122 ( BL122, BLN122, WL62);
sram_cell_6t_3 inst_cell_62_121 ( BL121, BLN121, WL62);
sram_cell_6t_3 inst_cell_62_120 ( BL120, BLN120, WL62);
sram_cell_6t_3 inst_cell_62_119 ( BL119, BLN119, WL62);
sram_cell_6t_3 inst_cell_62_118 ( BL118, BLN118, WL62);
sram_cell_6t_3 inst_cell_62_117 ( BL117, BLN117, WL62);
sram_cell_6t_3 inst_cell_62_116 ( BL116, BLN116, WL62);
sram_cell_6t_3 inst_cell_62_115 ( BL115, BLN115, WL62);
sram_cell_6t_3 inst_cell_62_114 ( BL114, BLN114, WL62);
sram_cell_6t_3 inst_cell_62_113 ( BL113, BLN113, WL62);
sram_cell_6t_3 inst_cell_62_112 ( BL112, BLN112, WL62);
sram_cell_6t_3 inst_cell_62_111 ( BL111, BLN111, WL62);
sram_cell_6t_3 inst_cell_62_110 ( BL110, BLN110, WL62);
sram_cell_6t_3 inst_cell_62_109 ( BL109, BLN109, WL62);
sram_cell_6t_3 inst_cell_62_108 ( BL108, BLN108, WL62);
sram_cell_6t_3 inst_cell_62_107 ( BL107, BLN107, WL62);
sram_cell_6t_3 inst_cell_62_106 ( BL106, BLN106, WL62);
sram_cell_6t_3 inst_cell_62_105 ( BL105, BLN105, WL62);
sram_cell_6t_3 inst_cell_62_104 ( BL104, BLN104, WL62);
sram_cell_6t_3 inst_cell_62_103 ( BL103, BLN103, WL62);
sram_cell_6t_3 inst_cell_62_102 ( BL102, BLN102, WL62);
sram_cell_6t_3 inst_cell_62_101 ( BL101, BLN101, WL62);
sram_cell_6t_3 inst_cell_62_100 ( BL100, BLN100, WL62);
sram_cell_6t_3 inst_cell_62_99 ( BL99, BLN99, WL62);
sram_cell_6t_3 inst_cell_62_98 ( BL98, BLN98, WL62);
sram_cell_6t_3 inst_cell_62_97 ( BL97, BLN97, WL62);
sram_cell_6t_3 inst_cell_62_96 ( BL96, BLN96, WL62);
sram_cell_6t_3 inst_cell_62_95 ( BL95, BLN95, WL62);
sram_cell_6t_3 inst_cell_62_94 ( BL94, BLN94, WL62);
sram_cell_6t_3 inst_cell_62_93 ( BL93, BLN93, WL62);
sram_cell_6t_3 inst_cell_62_92 ( BL92, BLN92, WL62);
sram_cell_6t_3 inst_cell_62_91 ( BL91, BLN91, WL62);
sram_cell_6t_3 inst_cell_62_90 ( BL90, BLN90, WL62);
sram_cell_6t_3 inst_cell_62_89 ( BL89, BLN89, WL62);
sram_cell_6t_3 inst_cell_62_88 ( BL88, BLN88, WL62);
sram_cell_6t_3 inst_cell_62_87 ( BL87, BLN87, WL62);
sram_cell_6t_3 inst_cell_62_86 ( BL86, BLN86, WL62);
sram_cell_6t_3 inst_cell_62_85 ( BL85, BLN85, WL62);
sram_cell_6t_3 inst_cell_62_84 ( BL84, BLN84, WL62);
sram_cell_6t_3 inst_cell_62_83 ( BL83, BLN83, WL62);
sram_cell_6t_3 inst_cell_62_82 ( BL82, BLN82, WL62);
sram_cell_6t_3 inst_cell_62_81 ( BL81, BLN81, WL62);
sram_cell_6t_3 inst_cell_62_80 ( BL80, BLN80, WL62);
sram_cell_6t_3 inst_cell_62_79 ( BL79, BLN79, WL62);
sram_cell_6t_3 inst_cell_62_78 ( BL78, BLN78, WL62);
sram_cell_6t_3 inst_cell_62_77 ( BL77, BLN77, WL62);
sram_cell_6t_3 inst_cell_62_76 ( BL76, BLN76, WL62);
sram_cell_6t_3 inst_cell_62_75 ( BL75, BLN75, WL62);
sram_cell_6t_3 inst_cell_62_74 ( BL74, BLN74, WL62);
sram_cell_6t_3 inst_cell_62_73 ( BL73, BLN73, WL62);
sram_cell_6t_3 inst_cell_62_72 ( BL72, BLN72, WL62);
sram_cell_6t_3 inst_cell_62_71 ( BL71, BLN71, WL62);
sram_cell_6t_3 inst_cell_62_70 ( BL70, BLN70, WL62);
sram_cell_6t_3 inst_cell_62_69 ( BL69, BLN69, WL62);
sram_cell_6t_3 inst_cell_62_68 ( BL68, BLN68, WL62);
sram_cell_6t_3 inst_cell_62_67 ( BL67, BLN67, WL62);
sram_cell_6t_3 inst_cell_62_66 ( BL66, BLN66, WL62);
sram_cell_6t_3 inst_cell_62_65 ( BL65, BLN65, WL62);
sram_cell_6t_3 inst_cell_62_64 ( BL64, BLN64, WL62);
sram_cell_6t_3 inst_cell_62_63 ( BL63, BLN63, WL62);
sram_cell_6t_3 inst_cell_62_62 ( BL62, BLN62, WL62);
sram_cell_6t_3 inst_cell_62_61 ( BL61, BLN61, WL62);
sram_cell_6t_3 inst_cell_62_60 ( BL60, BLN60, WL62);
sram_cell_6t_3 inst_cell_62_59 ( BL59, BLN59, WL62);
sram_cell_6t_3 inst_cell_62_58 ( BL58, BLN58, WL62);
sram_cell_6t_3 inst_cell_62_57 ( BL57, BLN57, WL62);
sram_cell_6t_3 inst_cell_62_56 ( BL56, BLN56, WL62);
sram_cell_6t_3 inst_cell_62_55 ( BL55, BLN55, WL62);
sram_cell_6t_3 inst_cell_62_54 ( BL54, BLN54, WL62);
sram_cell_6t_3 inst_cell_62_53 ( BL53, BLN53, WL62);
sram_cell_6t_3 inst_cell_62_52 ( BL52, BLN52, WL62);
sram_cell_6t_3 inst_cell_62_51 ( BL51, BLN51, WL62);
sram_cell_6t_3 inst_cell_62_50 ( BL50, BLN50, WL62);
sram_cell_6t_3 inst_cell_62_49 ( BL49, BLN49, WL62);
sram_cell_6t_3 inst_cell_62_48 ( BL48, BLN48, WL62);
sram_cell_6t_3 inst_cell_62_47 ( BL47, BLN47, WL62);
sram_cell_6t_3 inst_cell_62_46 ( BL46, BLN46, WL62);
sram_cell_6t_3 inst_cell_62_45 ( BL45, BLN45, WL62);
sram_cell_6t_3 inst_cell_62_44 ( BL44, BLN44, WL62);
sram_cell_6t_3 inst_cell_62_43 ( BL43, BLN43, WL62);
sram_cell_6t_3 inst_cell_62_42 ( BL42, BLN42, WL62);
sram_cell_6t_3 inst_cell_62_41 ( BL41, BLN41, WL62);
sram_cell_6t_3 inst_cell_62_40 ( BL40, BLN40, WL62);
sram_cell_6t_3 inst_cell_62_39 ( BL39, BLN39, WL62);
sram_cell_6t_3 inst_cell_62_38 ( BL38, BLN38, WL62);
sram_cell_6t_3 inst_cell_62_37 ( BL37, BLN37, WL62);
sram_cell_6t_3 inst_cell_62_36 ( BL36, BLN36, WL62);
sram_cell_6t_3 inst_cell_62_35 ( BL35, BLN35, WL62);
sram_cell_6t_3 inst_cell_62_34 ( BL34, BLN34, WL62);
sram_cell_6t_3 inst_cell_62_33 ( BL33, BLN33, WL62);
sram_cell_6t_3 inst_cell_62_32 ( BL32, BLN32, WL62);
sram_cell_6t_3 inst_cell_62_31 ( BL31, BLN31, WL62);
sram_cell_6t_3 inst_cell_62_30 ( BL30, BLN30, WL62);
sram_cell_6t_3 inst_cell_62_29 ( BL29, BLN29, WL62);
sram_cell_6t_3 inst_cell_62_28 ( BL28, BLN28, WL62);
sram_cell_6t_3 inst_cell_62_27 ( BL27, BLN27, WL62);
sram_cell_6t_3 inst_cell_62_26 ( BL26, BLN26, WL62);
sram_cell_6t_3 inst_cell_62_25 ( BL25, BLN25, WL62);
sram_cell_6t_3 inst_cell_62_24 ( BL24, BLN24, WL62);
sram_cell_6t_3 inst_cell_62_23 ( BL23, BLN23, WL62);
sram_cell_6t_3 inst_cell_62_22 ( BL22, BLN22, WL62);
sram_cell_6t_3 inst_cell_62_21 ( BL21, BLN21, WL62);
sram_cell_6t_3 inst_cell_62_20 ( BL20, BLN20, WL62);
sram_cell_6t_3 inst_cell_62_19 ( BL19, BLN19, WL62);
sram_cell_6t_3 inst_cell_62_18 ( BL18, BLN18, WL62);
sram_cell_6t_3 inst_cell_62_17 ( BL17, BLN17, WL62);
sram_cell_6t_3 inst_cell_62_16 ( BL16, BLN16, WL62);
sram_cell_6t_3 inst_cell_62_15 ( BL15, BLN15, WL62);
sram_cell_6t_3 inst_cell_62_14 ( BL14, BLN14, WL62);
sram_cell_6t_3 inst_cell_62_13 ( BL13, BLN13, WL62);
sram_cell_6t_3 inst_cell_62_12 ( BL12, BLN12, WL62);
sram_cell_6t_3 inst_cell_62_11 ( BL11, BLN11, WL62);
sram_cell_6t_3 inst_cell_62_10 ( BL10, BLN10, WL62);
sram_cell_6t_3 inst_cell_62_9 ( BL9, BLN9, WL62);
sram_cell_6t_3 inst_cell_62_8 ( BL8, BLN8, WL62);
sram_cell_6t_3 inst_cell_62_7 ( BL7, BLN7, WL62);
sram_cell_6t_3 inst_cell_62_6 ( BL6, BLN6, WL62);
sram_cell_6t_3 inst_cell_62_5 ( BL5, BLN5, WL62);
sram_cell_6t_3 inst_cell_62_4 ( BL4, BLN4, WL62);
sram_cell_6t_3 inst_cell_62_3 ( BL3, BLN3, WL62);
sram_cell_6t_3 inst_cell_62_2 ( BL2, BLN2, WL62);
sram_cell_6t_3 inst_cell_62_1 ( BL1, BLN1, WL62);
sram_cell_6t_3 inst_cell_62_0 ( BL0, BLN0, WL62);
sram_cell_6t_3 inst_cell_61_127 ( BL127, BLN127, WL61);
sram_cell_6t_3 inst_cell_61_126 ( BL126, BLN126, WL61);
sram_cell_6t_3 inst_cell_61_125 ( BL125, BLN125, WL61);
sram_cell_6t_3 inst_cell_61_124 ( BL124, BLN124, WL61);
sram_cell_6t_3 inst_cell_61_123 ( BL123, BLN123, WL61);
sram_cell_6t_3 inst_cell_61_122 ( BL122, BLN122, WL61);
sram_cell_6t_3 inst_cell_61_121 ( BL121, BLN121, WL61);
sram_cell_6t_3 inst_cell_61_120 ( BL120, BLN120, WL61);
sram_cell_6t_3 inst_cell_61_119 ( BL119, BLN119, WL61);
sram_cell_6t_3 inst_cell_61_118 ( BL118, BLN118, WL61);
sram_cell_6t_3 inst_cell_61_117 ( BL117, BLN117, WL61);
sram_cell_6t_3 inst_cell_61_116 ( BL116, BLN116, WL61);
sram_cell_6t_3 inst_cell_61_115 ( BL115, BLN115, WL61);
sram_cell_6t_3 inst_cell_61_114 ( BL114, BLN114, WL61);
sram_cell_6t_3 inst_cell_61_113 ( BL113, BLN113, WL61);
sram_cell_6t_3 inst_cell_61_112 ( BL112, BLN112, WL61);
sram_cell_6t_3 inst_cell_61_111 ( BL111, BLN111, WL61);
sram_cell_6t_3 inst_cell_61_110 ( BL110, BLN110, WL61);
sram_cell_6t_3 inst_cell_61_109 ( BL109, BLN109, WL61);
sram_cell_6t_3 inst_cell_61_108 ( BL108, BLN108, WL61);
sram_cell_6t_3 inst_cell_61_107 ( BL107, BLN107, WL61);
sram_cell_6t_3 inst_cell_61_106 ( BL106, BLN106, WL61);
sram_cell_6t_3 inst_cell_61_105 ( BL105, BLN105, WL61);
sram_cell_6t_3 inst_cell_61_104 ( BL104, BLN104, WL61);
sram_cell_6t_3 inst_cell_61_103 ( BL103, BLN103, WL61);
sram_cell_6t_3 inst_cell_61_102 ( BL102, BLN102, WL61);
sram_cell_6t_3 inst_cell_61_101 ( BL101, BLN101, WL61);
sram_cell_6t_3 inst_cell_61_100 ( BL100, BLN100, WL61);
sram_cell_6t_3 inst_cell_61_99 ( BL99, BLN99, WL61);
sram_cell_6t_3 inst_cell_61_98 ( BL98, BLN98, WL61);
sram_cell_6t_3 inst_cell_61_97 ( BL97, BLN97, WL61);
sram_cell_6t_3 inst_cell_61_96 ( BL96, BLN96, WL61);
sram_cell_6t_3 inst_cell_61_95 ( BL95, BLN95, WL61);
sram_cell_6t_3 inst_cell_61_94 ( BL94, BLN94, WL61);
sram_cell_6t_3 inst_cell_61_93 ( BL93, BLN93, WL61);
sram_cell_6t_3 inst_cell_61_92 ( BL92, BLN92, WL61);
sram_cell_6t_3 inst_cell_61_91 ( BL91, BLN91, WL61);
sram_cell_6t_3 inst_cell_61_90 ( BL90, BLN90, WL61);
sram_cell_6t_3 inst_cell_61_89 ( BL89, BLN89, WL61);
sram_cell_6t_3 inst_cell_61_88 ( BL88, BLN88, WL61);
sram_cell_6t_3 inst_cell_61_87 ( BL87, BLN87, WL61);
sram_cell_6t_3 inst_cell_61_86 ( BL86, BLN86, WL61);
sram_cell_6t_3 inst_cell_61_85 ( BL85, BLN85, WL61);
sram_cell_6t_3 inst_cell_61_84 ( BL84, BLN84, WL61);
sram_cell_6t_3 inst_cell_61_83 ( BL83, BLN83, WL61);
sram_cell_6t_3 inst_cell_61_82 ( BL82, BLN82, WL61);
sram_cell_6t_3 inst_cell_61_81 ( BL81, BLN81, WL61);
sram_cell_6t_3 inst_cell_61_80 ( BL80, BLN80, WL61);
sram_cell_6t_3 inst_cell_61_79 ( BL79, BLN79, WL61);
sram_cell_6t_3 inst_cell_61_78 ( BL78, BLN78, WL61);
sram_cell_6t_3 inst_cell_61_77 ( BL77, BLN77, WL61);
sram_cell_6t_3 inst_cell_61_76 ( BL76, BLN76, WL61);
sram_cell_6t_3 inst_cell_61_75 ( BL75, BLN75, WL61);
sram_cell_6t_3 inst_cell_61_74 ( BL74, BLN74, WL61);
sram_cell_6t_3 inst_cell_61_73 ( BL73, BLN73, WL61);
sram_cell_6t_3 inst_cell_61_72 ( BL72, BLN72, WL61);
sram_cell_6t_3 inst_cell_61_71 ( BL71, BLN71, WL61);
sram_cell_6t_3 inst_cell_61_70 ( BL70, BLN70, WL61);
sram_cell_6t_3 inst_cell_61_69 ( BL69, BLN69, WL61);
sram_cell_6t_3 inst_cell_61_68 ( BL68, BLN68, WL61);
sram_cell_6t_3 inst_cell_61_67 ( BL67, BLN67, WL61);
sram_cell_6t_3 inst_cell_61_66 ( BL66, BLN66, WL61);
sram_cell_6t_3 inst_cell_61_65 ( BL65, BLN65, WL61);
sram_cell_6t_3 inst_cell_61_64 ( BL64, BLN64, WL61);
sram_cell_6t_3 inst_cell_61_63 ( BL63, BLN63, WL61);
sram_cell_6t_3 inst_cell_61_62 ( BL62, BLN62, WL61);
sram_cell_6t_3 inst_cell_61_61 ( BL61, BLN61, WL61);
sram_cell_6t_3 inst_cell_61_60 ( BL60, BLN60, WL61);
sram_cell_6t_3 inst_cell_61_59 ( BL59, BLN59, WL61);
sram_cell_6t_3 inst_cell_61_58 ( BL58, BLN58, WL61);
sram_cell_6t_3 inst_cell_61_57 ( BL57, BLN57, WL61);
sram_cell_6t_3 inst_cell_61_56 ( BL56, BLN56, WL61);
sram_cell_6t_3 inst_cell_61_55 ( BL55, BLN55, WL61);
sram_cell_6t_3 inst_cell_61_54 ( BL54, BLN54, WL61);
sram_cell_6t_3 inst_cell_61_53 ( BL53, BLN53, WL61);
sram_cell_6t_3 inst_cell_61_52 ( BL52, BLN52, WL61);
sram_cell_6t_3 inst_cell_61_51 ( BL51, BLN51, WL61);
sram_cell_6t_3 inst_cell_61_50 ( BL50, BLN50, WL61);
sram_cell_6t_3 inst_cell_61_49 ( BL49, BLN49, WL61);
sram_cell_6t_3 inst_cell_61_48 ( BL48, BLN48, WL61);
sram_cell_6t_3 inst_cell_61_47 ( BL47, BLN47, WL61);
sram_cell_6t_3 inst_cell_61_46 ( BL46, BLN46, WL61);
sram_cell_6t_3 inst_cell_61_45 ( BL45, BLN45, WL61);
sram_cell_6t_3 inst_cell_61_44 ( BL44, BLN44, WL61);
sram_cell_6t_3 inst_cell_61_43 ( BL43, BLN43, WL61);
sram_cell_6t_3 inst_cell_61_42 ( BL42, BLN42, WL61);
sram_cell_6t_3 inst_cell_61_41 ( BL41, BLN41, WL61);
sram_cell_6t_3 inst_cell_61_40 ( BL40, BLN40, WL61);
sram_cell_6t_3 inst_cell_61_39 ( BL39, BLN39, WL61);
sram_cell_6t_3 inst_cell_61_38 ( BL38, BLN38, WL61);
sram_cell_6t_3 inst_cell_61_37 ( BL37, BLN37, WL61);
sram_cell_6t_3 inst_cell_61_36 ( BL36, BLN36, WL61);
sram_cell_6t_3 inst_cell_61_35 ( BL35, BLN35, WL61);
sram_cell_6t_3 inst_cell_61_34 ( BL34, BLN34, WL61);
sram_cell_6t_3 inst_cell_61_33 ( BL33, BLN33, WL61);
sram_cell_6t_3 inst_cell_61_32 ( BL32, BLN32, WL61);
sram_cell_6t_3 inst_cell_61_31 ( BL31, BLN31, WL61);
sram_cell_6t_3 inst_cell_61_30 ( BL30, BLN30, WL61);
sram_cell_6t_3 inst_cell_61_29 ( BL29, BLN29, WL61);
sram_cell_6t_3 inst_cell_61_28 ( BL28, BLN28, WL61);
sram_cell_6t_3 inst_cell_61_27 ( BL27, BLN27, WL61);
sram_cell_6t_3 inst_cell_61_26 ( BL26, BLN26, WL61);
sram_cell_6t_3 inst_cell_61_25 ( BL25, BLN25, WL61);
sram_cell_6t_3 inst_cell_61_24 ( BL24, BLN24, WL61);
sram_cell_6t_3 inst_cell_61_23 ( BL23, BLN23, WL61);
sram_cell_6t_3 inst_cell_61_22 ( BL22, BLN22, WL61);
sram_cell_6t_3 inst_cell_61_21 ( BL21, BLN21, WL61);
sram_cell_6t_3 inst_cell_61_20 ( BL20, BLN20, WL61);
sram_cell_6t_3 inst_cell_61_19 ( BL19, BLN19, WL61);
sram_cell_6t_3 inst_cell_61_18 ( BL18, BLN18, WL61);
sram_cell_6t_3 inst_cell_61_17 ( BL17, BLN17, WL61);
sram_cell_6t_3 inst_cell_61_16 ( BL16, BLN16, WL61);
sram_cell_6t_3 inst_cell_61_15 ( BL15, BLN15, WL61);
sram_cell_6t_3 inst_cell_61_14 ( BL14, BLN14, WL61);
sram_cell_6t_3 inst_cell_61_13 ( BL13, BLN13, WL61);
sram_cell_6t_3 inst_cell_61_12 ( BL12, BLN12, WL61);
sram_cell_6t_3 inst_cell_61_11 ( BL11, BLN11, WL61);
sram_cell_6t_3 inst_cell_61_10 ( BL10, BLN10, WL61);
sram_cell_6t_3 inst_cell_61_9 ( BL9, BLN9, WL61);
sram_cell_6t_3 inst_cell_61_8 ( BL8, BLN8, WL61);
sram_cell_6t_3 inst_cell_61_7 ( BL7, BLN7, WL61);
sram_cell_6t_3 inst_cell_61_6 ( BL6, BLN6, WL61);
sram_cell_6t_3 inst_cell_61_5 ( BL5, BLN5, WL61);
sram_cell_6t_3 inst_cell_61_4 ( BL4, BLN4, WL61);
sram_cell_6t_3 inst_cell_61_3 ( BL3, BLN3, WL61);
sram_cell_6t_3 inst_cell_61_2 ( BL2, BLN2, WL61);
sram_cell_6t_3 inst_cell_61_1 ( BL1, BLN1, WL61);
sram_cell_6t_3 inst_cell_61_0 ( BL0, BLN0, WL61);
sram_cell_6t_3 inst_cell_60_127 ( BL127, BLN127, WL60);
sram_cell_6t_3 inst_cell_60_126 ( BL126, BLN126, WL60);
sram_cell_6t_3 inst_cell_60_125 ( BL125, BLN125, WL60);
sram_cell_6t_3 inst_cell_60_124 ( BL124, BLN124, WL60);
sram_cell_6t_3 inst_cell_60_123 ( BL123, BLN123, WL60);
sram_cell_6t_3 inst_cell_60_122 ( BL122, BLN122, WL60);
sram_cell_6t_3 inst_cell_60_121 ( BL121, BLN121, WL60);
sram_cell_6t_3 inst_cell_60_120 ( BL120, BLN120, WL60);
sram_cell_6t_3 inst_cell_60_119 ( BL119, BLN119, WL60);
sram_cell_6t_3 inst_cell_60_118 ( BL118, BLN118, WL60);
sram_cell_6t_3 inst_cell_60_117 ( BL117, BLN117, WL60);
sram_cell_6t_3 inst_cell_60_116 ( BL116, BLN116, WL60);
sram_cell_6t_3 inst_cell_60_115 ( BL115, BLN115, WL60);
sram_cell_6t_3 inst_cell_60_114 ( BL114, BLN114, WL60);
sram_cell_6t_3 inst_cell_60_113 ( BL113, BLN113, WL60);
sram_cell_6t_3 inst_cell_60_112 ( BL112, BLN112, WL60);
sram_cell_6t_3 inst_cell_60_111 ( BL111, BLN111, WL60);
sram_cell_6t_3 inst_cell_60_110 ( BL110, BLN110, WL60);
sram_cell_6t_3 inst_cell_60_109 ( BL109, BLN109, WL60);
sram_cell_6t_3 inst_cell_60_108 ( BL108, BLN108, WL60);
sram_cell_6t_3 inst_cell_60_107 ( BL107, BLN107, WL60);
sram_cell_6t_3 inst_cell_60_106 ( BL106, BLN106, WL60);
sram_cell_6t_3 inst_cell_60_105 ( BL105, BLN105, WL60);
sram_cell_6t_3 inst_cell_60_104 ( BL104, BLN104, WL60);
sram_cell_6t_3 inst_cell_60_103 ( BL103, BLN103, WL60);
sram_cell_6t_3 inst_cell_60_102 ( BL102, BLN102, WL60);
sram_cell_6t_3 inst_cell_60_101 ( BL101, BLN101, WL60);
sram_cell_6t_3 inst_cell_60_100 ( BL100, BLN100, WL60);
sram_cell_6t_3 inst_cell_60_99 ( BL99, BLN99, WL60);
sram_cell_6t_3 inst_cell_60_98 ( BL98, BLN98, WL60);
sram_cell_6t_3 inst_cell_60_97 ( BL97, BLN97, WL60);
sram_cell_6t_3 inst_cell_60_96 ( BL96, BLN96, WL60);
sram_cell_6t_3 inst_cell_60_95 ( BL95, BLN95, WL60);
sram_cell_6t_3 inst_cell_60_94 ( BL94, BLN94, WL60);
sram_cell_6t_3 inst_cell_60_93 ( BL93, BLN93, WL60);
sram_cell_6t_3 inst_cell_60_92 ( BL92, BLN92, WL60);
sram_cell_6t_3 inst_cell_60_91 ( BL91, BLN91, WL60);
sram_cell_6t_3 inst_cell_60_90 ( BL90, BLN90, WL60);
sram_cell_6t_3 inst_cell_60_89 ( BL89, BLN89, WL60);
sram_cell_6t_3 inst_cell_60_88 ( BL88, BLN88, WL60);
sram_cell_6t_3 inst_cell_60_87 ( BL87, BLN87, WL60);
sram_cell_6t_3 inst_cell_60_86 ( BL86, BLN86, WL60);
sram_cell_6t_3 inst_cell_60_85 ( BL85, BLN85, WL60);
sram_cell_6t_3 inst_cell_60_84 ( BL84, BLN84, WL60);
sram_cell_6t_3 inst_cell_60_83 ( BL83, BLN83, WL60);
sram_cell_6t_3 inst_cell_60_82 ( BL82, BLN82, WL60);
sram_cell_6t_3 inst_cell_60_81 ( BL81, BLN81, WL60);
sram_cell_6t_3 inst_cell_60_80 ( BL80, BLN80, WL60);
sram_cell_6t_3 inst_cell_60_79 ( BL79, BLN79, WL60);
sram_cell_6t_3 inst_cell_60_78 ( BL78, BLN78, WL60);
sram_cell_6t_3 inst_cell_60_77 ( BL77, BLN77, WL60);
sram_cell_6t_3 inst_cell_60_76 ( BL76, BLN76, WL60);
sram_cell_6t_3 inst_cell_60_75 ( BL75, BLN75, WL60);
sram_cell_6t_3 inst_cell_60_74 ( BL74, BLN74, WL60);
sram_cell_6t_3 inst_cell_60_73 ( BL73, BLN73, WL60);
sram_cell_6t_3 inst_cell_60_72 ( BL72, BLN72, WL60);
sram_cell_6t_3 inst_cell_60_71 ( BL71, BLN71, WL60);
sram_cell_6t_3 inst_cell_60_70 ( BL70, BLN70, WL60);
sram_cell_6t_3 inst_cell_60_69 ( BL69, BLN69, WL60);
sram_cell_6t_3 inst_cell_60_68 ( BL68, BLN68, WL60);
sram_cell_6t_3 inst_cell_60_67 ( BL67, BLN67, WL60);
sram_cell_6t_3 inst_cell_60_66 ( BL66, BLN66, WL60);
sram_cell_6t_3 inst_cell_60_65 ( BL65, BLN65, WL60);
sram_cell_6t_3 inst_cell_60_64 ( BL64, BLN64, WL60);
sram_cell_6t_3 inst_cell_60_63 ( BL63, BLN63, WL60);
sram_cell_6t_3 inst_cell_60_62 ( BL62, BLN62, WL60);
sram_cell_6t_3 inst_cell_60_61 ( BL61, BLN61, WL60);
sram_cell_6t_3 inst_cell_60_60 ( BL60, BLN60, WL60);
sram_cell_6t_3 inst_cell_60_59 ( BL59, BLN59, WL60);
sram_cell_6t_3 inst_cell_60_58 ( BL58, BLN58, WL60);
sram_cell_6t_3 inst_cell_60_57 ( BL57, BLN57, WL60);
sram_cell_6t_3 inst_cell_60_56 ( BL56, BLN56, WL60);
sram_cell_6t_3 inst_cell_60_55 ( BL55, BLN55, WL60);
sram_cell_6t_3 inst_cell_60_54 ( BL54, BLN54, WL60);
sram_cell_6t_3 inst_cell_60_53 ( BL53, BLN53, WL60);
sram_cell_6t_3 inst_cell_60_52 ( BL52, BLN52, WL60);
sram_cell_6t_3 inst_cell_60_51 ( BL51, BLN51, WL60);
sram_cell_6t_3 inst_cell_60_50 ( BL50, BLN50, WL60);
sram_cell_6t_3 inst_cell_60_49 ( BL49, BLN49, WL60);
sram_cell_6t_3 inst_cell_60_48 ( BL48, BLN48, WL60);
sram_cell_6t_3 inst_cell_60_47 ( BL47, BLN47, WL60);
sram_cell_6t_3 inst_cell_60_46 ( BL46, BLN46, WL60);
sram_cell_6t_3 inst_cell_60_45 ( BL45, BLN45, WL60);
sram_cell_6t_3 inst_cell_60_44 ( BL44, BLN44, WL60);
sram_cell_6t_3 inst_cell_60_43 ( BL43, BLN43, WL60);
sram_cell_6t_3 inst_cell_60_42 ( BL42, BLN42, WL60);
sram_cell_6t_3 inst_cell_60_41 ( BL41, BLN41, WL60);
sram_cell_6t_3 inst_cell_60_40 ( BL40, BLN40, WL60);
sram_cell_6t_3 inst_cell_60_39 ( BL39, BLN39, WL60);
sram_cell_6t_3 inst_cell_60_38 ( BL38, BLN38, WL60);
sram_cell_6t_3 inst_cell_60_37 ( BL37, BLN37, WL60);
sram_cell_6t_3 inst_cell_60_36 ( BL36, BLN36, WL60);
sram_cell_6t_3 inst_cell_60_35 ( BL35, BLN35, WL60);
sram_cell_6t_3 inst_cell_60_34 ( BL34, BLN34, WL60);
sram_cell_6t_3 inst_cell_60_33 ( BL33, BLN33, WL60);
sram_cell_6t_3 inst_cell_60_32 ( BL32, BLN32, WL60);
sram_cell_6t_3 inst_cell_60_31 ( BL31, BLN31, WL60);
sram_cell_6t_3 inst_cell_60_30 ( BL30, BLN30, WL60);
sram_cell_6t_3 inst_cell_60_29 ( BL29, BLN29, WL60);
sram_cell_6t_3 inst_cell_60_28 ( BL28, BLN28, WL60);
sram_cell_6t_3 inst_cell_60_27 ( BL27, BLN27, WL60);
sram_cell_6t_3 inst_cell_60_26 ( BL26, BLN26, WL60);
sram_cell_6t_3 inst_cell_60_25 ( BL25, BLN25, WL60);
sram_cell_6t_3 inst_cell_60_24 ( BL24, BLN24, WL60);
sram_cell_6t_3 inst_cell_60_23 ( BL23, BLN23, WL60);
sram_cell_6t_3 inst_cell_60_22 ( BL22, BLN22, WL60);
sram_cell_6t_3 inst_cell_60_21 ( BL21, BLN21, WL60);
sram_cell_6t_3 inst_cell_60_20 ( BL20, BLN20, WL60);
sram_cell_6t_3 inst_cell_60_19 ( BL19, BLN19, WL60);
sram_cell_6t_3 inst_cell_60_18 ( BL18, BLN18, WL60);
sram_cell_6t_3 inst_cell_60_17 ( BL17, BLN17, WL60);
sram_cell_6t_3 inst_cell_60_16 ( BL16, BLN16, WL60);
sram_cell_6t_3 inst_cell_60_15 ( BL15, BLN15, WL60);
sram_cell_6t_3 inst_cell_60_14 ( BL14, BLN14, WL60);
sram_cell_6t_3 inst_cell_60_13 ( BL13, BLN13, WL60);
sram_cell_6t_3 inst_cell_60_12 ( BL12, BLN12, WL60);
sram_cell_6t_3 inst_cell_60_11 ( BL11, BLN11, WL60);
sram_cell_6t_3 inst_cell_60_10 ( BL10, BLN10, WL60);
sram_cell_6t_3 inst_cell_60_9 ( BL9, BLN9, WL60);
sram_cell_6t_3 inst_cell_60_8 ( BL8, BLN8, WL60);
sram_cell_6t_3 inst_cell_60_7 ( BL7, BLN7, WL60);
sram_cell_6t_3 inst_cell_60_6 ( BL6, BLN6, WL60);
sram_cell_6t_3 inst_cell_60_5 ( BL5, BLN5, WL60);
sram_cell_6t_3 inst_cell_60_4 ( BL4, BLN4, WL60);
sram_cell_6t_3 inst_cell_60_3 ( BL3, BLN3, WL60);
sram_cell_6t_3 inst_cell_60_2 ( BL2, BLN2, WL60);
sram_cell_6t_3 inst_cell_60_1 ( BL1, BLN1, WL60);
sram_cell_6t_3 inst_cell_60_0 ( BL0, BLN0, WL60);
sram_cell_6t_3 inst_cell_59_127 ( BL127, BLN127, WL59);
sram_cell_6t_3 inst_cell_59_126 ( BL126, BLN126, WL59);
sram_cell_6t_3 inst_cell_59_125 ( BL125, BLN125, WL59);
sram_cell_6t_3 inst_cell_59_124 ( BL124, BLN124, WL59);
sram_cell_6t_3 inst_cell_59_123 ( BL123, BLN123, WL59);
sram_cell_6t_3 inst_cell_59_122 ( BL122, BLN122, WL59);
sram_cell_6t_3 inst_cell_59_121 ( BL121, BLN121, WL59);
sram_cell_6t_3 inst_cell_59_120 ( BL120, BLN120, WL59);
sram_cell_6t_3 inst_cell_59_119 ( BL119, BLN119, WL59);
sram_cell_6t_3 inst_cell_59_118 ( BL118, BLN118, WL59);
sram_cell_6t_3 inst_cell_59_117 ( BL117, BLN117, WL59);
sram_cell_6t_3 inst_cell_59_116 ( BL116, BLN116, WL59);
sram_cell_6t_3 inst_cell_59_115 ( BL115, BLN115, WL59);
sram_cell_6t_3 inst_cell_59_114 ( BL114, BLN114, WL59);
sram_cell_6t_3 inst_cell_59_113 ( BL113, BLN113, WL59);
sram_cell_6t_3 inst_cell_59_112 ( BL112, BLN112, WL59);
sram_cell_6t_3 inst_cell_59_111 ( BL111, BLN111, WL59);
sram_cell_6t_3 inst_cell_59_110 ( BL110, BLN110, WL59);
sram_cell_6t_3 inst_cell_59_109 ( BL109, BLN109, WL59);
sram_cell_6t_3 inst_cell_59_108 ( BL108, BLN108, WL59);
sram_cell_6t_3 inst_cell_59_107 ( BL107, BLN107, WL59);
sram_cell_6t_3 inst_cell_59_106 ( BL106, BLN106, WL59);
sram_cell_6t_3 inst_cell_59_105 ( BL105, BLN105, WL59);
sram_cell_6t_3 inst_cell_59_104 ( BL104, BLN104, WL59);
sram_cell_6t_3 inst_cell_59_103 ( BL103, BLN103, WL59);
sram_cell_6t_3 inst_cell_59_102 ( BL102, BLN102, WL59);
sram_cell_6t_3 inst_cell_59_101 ( BL101, BLN101, WL59);
sram_cell_6t_3 inst_cell_59_100 ( BL100, BLN100, WL59);
sram_cell_6t_3 inst_cell_59_99 ( BL99, BLN99, WL59);
sram_cell_6t_3 inst_cell_59_98 ( BL98, BLN98, WL59);
sram_cell_6t_3 inst_cell_59_97 ( BL97, BLN97, WL59);
sram_cell_6t_3 inst_cell_59_96 ( BL96, BLN96, WL59);
sram_cell_6t_3 inst_cell_59_95 ( BL95, BLN95, WL59);
sram_cell_6t_3 inst_cell_59_94 ( BL94, BLN94, WL59);
sram_cell_6t_3 inst_cell_59_93 ( BL93, BLN93, WL59);
sram_cell_6t_3 inst_cell_59_92 ( BL92, BLN92, WL59);
sram_cell_6t_3 inst_cell_59_91 ( BL91, BLN91, WL59);
sram_cell_6t_3 inst_cell_59_90 ( BL90, BLN90, WL59);
sram_cell_6t_3 inst_cell_59_89 ( BL89, BLN89, WL59);
sram_cell_6t_3 inst_cell_59_88 ( BL88, BLN88, WL59);
sram_cell_6t_3 inst_cell_59_87 ( BL87, BLN87, WL59);
sram_cell_6t_3 inst_cell_59_86 ( BL86, BLN86, WL59);
sram_cell_6t_3 inst_cell_59_85 ( BL85, BLN85, WL59);
sram_cell_6t_3 inst_cell_59_84 ( BL84, BLN84, WL59);
sram_cell_6t_3 inst_cell_59_83 ( BL83, BLN83, WL59);
sram_cell_6t_3 inst_cell_59_82 ( BL82, BLN82, WL59);
sram_cell_6t_3 inst_cell_59_81 ( BL81, BLN81, WL59);
sram_cell_6t_3 inst_cell_59_80 ( BL80, BLN80, WL59);
sram_cell_6t_3 inst_cell_59_79 ( BL79, BLN79, WL59);
sram_cell_6t_3 inst_cell_59_78 ( BL78, BLN78, WL59);
sram_cell_6t_3 inst_cell_59_77 ( BL77, BLN77, WL59);
sram_cell_6t_3 inst_cell_59_76 ( BL76, BLN76, WL59);
sram_cell_6t_3 inst_cell_59_75 ( BL75, BLN75, WL59);
sram_cell_6t_3 inst_cell_59_74 ( BL74, BLN74, WL59);
sram_cell_6t_3 inst_cell_59_73 ( BL73, BLN73, WL59);
sram_cell_6t_3 inst_cell_59_72 ( BL72, BLN72, WL59);
sram_cell_6t_3 inst_cell_59_71 ( BL71, BLN71, WL59);
sram_cell_6t_3 inst_cell_59_70 ( BL70, BLN70, WL59);
sram_cell_6t_3 inst_cell_59_69 ( BL69, BLN69, WL59);
sram_cell_6t_3 inst_cell_59_68 ( BL68, BLN68, WL59);
sram_cell_6t_3 inst_cell_59_67 ( BL67, BLN67, WL59);
sram_cell_6t_3 inst_cell_59_66 ( BL66, BLN66, WL59);
sram_cell_6t_3 inst_cell_59_65 ( BL65, BLN65, WL59);
sram_cell_6t_3 inst_cell_59_64 ( BL64, BLN64, WL59);
sram_cell_6t_3 inst_cell_59_63 ( BL63, BLN63, WL59);
sram_cell_6t_3 inst_cell_59_62 ( BL62, BLN62, WL59);
sram_cell_6t_3 inst_cell_59_61 ( BL61, BLN61, WL59);
sram_cell_6t_3 inst_cell_59_60 ( BL60, BLN60, WL59);
sram_cell_6t_3 inst_cell_59_59 ( BL59, BLN59, WL59);
sram_cell_6t_3 inst_cell_59_58 ( BL58, BLN58, WL59);
sram_cell_6t_3 inst_cell_59_57 ( BL57, BLN57, WL59);
sram_cell_6t_3 inst_cell_59_56 ( BL56, BLN56, WL59);
sram_cell_6t_3 inst_cell_59_55 ( BL55, BLN55, WL59);
sram_cell_6t_3 inst_cell_59_54 ( BL54, BLN54, WL59);
sram_cell_6t_3 inst_cell_59_53 ( BL53, BLN53, WL59);
sram_cell_6t_3 inst_cell_59_52 ( BL52, BLN52, WL59);
sram_cell_6t_3 inst_cell_59_51 ( BL51, BLN51, WL59);
sram_cell_6t_3 inst_cell_59_50 ( BL50, BLN50, WL59);
sram_cell_6t_3 inst_cell_59_49 ( BL49, BLN49, WL59);
sram_cell_6t_3 inst_cell_59_48 ( BL48, BLN48, WL59);
sram_cell_6t_3 inst_cell_59_47 ( BL47, BLN47, WL59);
sram_cell_6t_3 inst_cell_59_46 ( BL46, BLN46, WL59);
sram_cell_6t_3 inst_cell_59_45 ( BL45, BLN45, WL59);
sram_cell_6t_3 inst_cell_59_44 ( BL44, BLN44, WL59);
sram_cell_6t_3 inst_cell_59_43 ( BL43, BLN43, WL59);
sram_cell_6t_3 inst_cell_59_42 ( BL42, BLN42, WL59);
sram_cell_6t_3 inst_cell_59_41 ( BL41, BLN41, WL59);
sram_cell_6t_3 inst_cell_59_40 ( BL40, BLN40, WL59);
sram_cell_6t_3 inst_cell_59_39 ( BL39, BLN39, WL59);
sram_cell_6t_3 inst_cell_59_38 ( BL38, BLN38, WL59);
sram_cell_6t_3 inst_cell_59_37 ( BL37, BLN37, WL59);
sram_cell_6t_3 inst_cell_59_36 ( BL36, BLN36, WL59);
sram_cell_6t_3 inst_cell_59_35 ( BL35, BLN35, WL59);
sram_cell_6t_3 inst_cell_59_34 ( BL34, BLN34, WL59);
sram_cell_6t_3 inst_cell_59_33 ( BL33, BLN33, WL59);
sram_cell_6t_3 inst_cell_59_32 ( BL32, BLN32, WL59);
sram_cell_6t_3 inst_cell_59_31 ( BL31, BLN31, WL59);
sram_cell_6t_3 inst_cell_59_30 ( BL30, BLN30, WL59);
sram_cell_6t_3 inst_cell_59_29 ( BL29, BLN29, WL59);
sram_cell_6t_3 inst_cell_59_28 ( BL28, BLN28, WL59);
sram_cell_6t_3 inst_cell_59_27 ( BL27, BLN27, WL59);
sram_cell_6t_3 inst_cell_59_26 ( BL26, BLN26, WL59);
sram_cell_6t_3 inst_cell_59_25 ( BL25, BLN25, WL59);
sram_cell_6t_3 inst_cell_59_24 ( BL24, BLN24, WL59);
sram_cell_6t_3 inst_cell_59_23 ( BL23, BLN23, WL59);
sram_cell_6t_3 inst_cell_59_22 ( BL22, BLN22, WL59);
sram_cell_6t_3 inst_cell_59_21 ( BL21, BLN21, WL59);
sram_cell_6t_3 inst_cell_59_20 ( BL20, BLN20, WL59);
sram_cell_6t_3 inst_cell_59_19 ( BL19, BLN19, WL59);
sram_cell_6t_3 inst_cell_59_18 ( BL18, BLN18, WL59);
sram_cell_6t_3 inst_cell_59_17 ( BL17, BLN17, WL59);
sram_cell_6t_3 inst_cell_59_16 ( BL16, BLN16, WL59);
sram_cell_6t_3 inst_cell_59_15 ( BL15, BLN15, WL59);
sram_cell_6t_3 inst_cell_59_14 ( BL14, BLN14, WL59);
sram_cell_6t_3 inst_cell_59_13 ( BL13, BLN13, WL59);
sram_cell_6t_3 inst_cell_59_12 ( BL12, BLN12, WL59);
sram_cell_6t_3 inst_cell_59_11 ( BL11, BLN11, WL59);
sram_cell_6t_3 inst_cell_59_10 ( BL10, BLN10, WL59);
sram_cell_6t_3 inst_cell_59_9 ( BL9, BLN9, WL59);
sram_cell_6t_3 inst_cell_59_8 ( BL8, BLN8, WL59);
sram_cell_6t_3 inst_cell_59_7 ( BL7, BLN7, WL59);
sram_cell_6t_3 inst_cell_59_6 ( BL6, BLN6, WL59);
sram_cell_6t_3 inst_cell_59_5 ( BL5, BLN5, WL59);
sram_cell_6t_3 inst_cell_59_4 ( BL4, BLN4, WL59);
sram_cell_6t_3 inst_cell_59_3 ( BL3, BLN3, WL59);
sram_cell_6t_3 inst_cell_59_2 ( BL2, BLN2, WL59);
sram_cell_6t_3 inst_cell_59_1 ( BL1, BLN1, WL59);
sram_cell_6t_3 inst_cell_59_0 ( BL0, BLN0, WL59);
sram_cell_6t_3 inst_cell_58_127 ( BL127, BLN127, WL58);
sram_cell_6t_3 inst_cell_58_126 ( BL126, BLN126, WL58);
sram_cell_6t_3 inst_cell_58_125 ( BL125, BLN125, WL58);
sram_cell_6t_3 inst_cell_58_124 ( BL124, BLN124, WL58);
sram_cell_6t_3 inst_cell_58_123 ( BL123, BLN123, WL58);
sram_cell_6t_3 inst_cell_58_122 ( BL122, BLN122, WL58);
sram_cell_6t_3 inst_cell_58_121 ( BL121, BLN121, WL58);
sram_cell_6t_3 inst_cell_58_120 ( BL120, BLN120, WL58);
sram_cell_6t_3 inst_cell_58_119 ( BL119, BLN119, WL58);
sram_cell_6t_3 inst_cell_58_118 ( BL118, BLN118, WL58);
sram_cell_6t_3 inst_cell_58_117 ( BL117, BLN117, WL58);
sram_cell_6t_3 inst_cell_58_116 ( BL116, BLN116, WL58);
sram_cell_6t_3 inst_cell_58_115 ( BL115, BLN115, WL58);
sram_cell_6t_3 inst_cell_58_114 ( BL114, BLN114, WL58);
sram_cell_6t_3 inst_cell_58_113 ( BL113, BLN113, WL58);
sram_cell_6t_3 inst_cell_58_112 ( BL112, BLN112, WL58);
sram_cell_6t_3 inst_cell_58_111 ( BL111, BLN111, WL58);
sram_cell_6t_3 inst_cell_58_110 ( BL110, BLN110, WL58);
sram_cell_6t_3 inst_cell_58_109 ( BL109, BLN109, WL58);
sram_cell_6t_3 inst_cell_58_108 ( BL108, BLN108, WL58);
sram_cell_6t_3 inst_cell_58_107 ( BL107, BLN107, WL58);
sram_cell_6t_3 inst_cell_58_106 ( BL106, BLN106, WL58);
sram_cell_6t_3 inst_cell_58_105 ( BL105, BLN105, WL58);
sram_cell_6t_3 inst_cell_58_104 ( BL104, BLN104, WL58);
sram_cell_6t_3 inst_cell_58_103 ( BL103, BLN103, WL58);
sram_cell_6t_3 inst_cell_58_102 ( BL102, BLN102, WL58);
sram_cell_6t_3 inst_cell_58_101 ( BL101, BLN101, WL58);
sram_cell_6t_3 inst_cell_58_100 ( BL100, BLN100, WL58);
sram_cell_6t_3 inst_cell_58_99 ( BL99, BLN99, WL58);
sram_cell_6t_3 inst_cell_58_98 ( BL98, BLN98, WL58);
sram_cell_6t_3 inst_cell_58_97 ( BL97, BLN97, WL58);
sram_cell_6t_3 inst_cell_58_96 ( BL96, BLN96, WL58);
sram_cell_6t_3 inst_cell_58_95 ( BL95, BLN95, WL58);
sram_cell_6t_3 inst_cell_58_94 ( BL94, BLN94, WL58);
sram_cell_6t_3 inst_cell_58_93 ( BL93, BLN93, WL58);
sram_cell_6t_3 inst_cell_58_92 ( BL92, BLN92, WL58);
sram_cell_6t_3 inst_cell_58_91 ( BL91, BLN91, WL58);
sram_cell_6t_3 inst_cell_58_90 ( BL90, BLN90, WL58);
sram_cell_6t_3 inst_cell_58_89 ( BL89, BLN89, WL58);
sram_cell_6t_3 inst_cell_58_88 ( BL88, BLN88, WL58);
sram_cell_6t_3 inst_cell_58_87 ( BL87, BLN87, WL58);
sram_cell_6t_3 inst_cell_58_86 ( BL86, BLN86, WL58);
sram_cell_6t_3 inst_cell_58_85 ( BL85, BLN85, WL58);
sram_cell_6t_3 inst_cell_58_84 ( BL84, BLN84, WL58);
sram_cell_6t_3 inst_cell_58_83 ( BL83, BLN83, WL58);
sram_cell_6t_3 inst_cell_58_82 ( BL82, BLN82, WL58);
sram_cell_6t_3 inst_cell_58_81 ( BL81, BLN81, WL58);
sram_cell_6t_3 inst_cell_58_80 ( BL80, BLN80, WL58);
sram_cell_6t_3 inst_cell_58_79 ( BL79, BLN79, WL58);
sram_cell_6t_3 inst_cell_58_78 ( BL78, BLN78, WL58);
sram_cell_6t_3 inst_cell_58_77 ( BL77, BLN77, WL58);
sram_cell_6t_3 inst_cell_58_76 ( BL76, BLN76, WL58);
sram_cell_6t_3 inst_cell_58_75 ( BL75, BLN75, WL58);
sram_cell_6t_3 inst_cell_58_74 ( BL74, BLN74, WL58);
sram_cell_6t_3 inst_cell_58_73 ( BL73, BLN73, WL58);
sram_cell_6t_3 inst_cell_58_72 ( BL72, BLN72, WL58);
sram_cell_6t_3 inst_cell_58_71 ( BL71, BLN71, WL58);
sram_cell_6t_3 inst_cell_58_70 ( BL70, BLN70, WL58);
sram_cell_6t_3 inst_cell_58_69 ( BL69, BLN69, WL58);
sram_cell_6t_3 inst_cell_58_68 ( BL68, BLN68, WL58);
sram_cell_6t_3 inst_cell_58_67 ( BL67, BLN67, WL58);
sram_cell_6t_3 inst_cell_58_66 ( BL66, BLN66, WL58);
sram_cell_6t_3 inst_cell_58_65 ( BL65, BLN65, WL58);
sram_cell_6t_3 inst_cell_58_64 ( BL64, BLN64, WL58);
sram_cell_6t_3 inst_cell_58_63 ( BL63, BLN63, WL58);
sram_cell_6t_3 inst_cell_58_62 ( BL62, BLN62, WL58);
sram_cell_6t_3 inst_cell_58_61 ( BL61, BLN61, WL58);
sram_cell_6t_3 inst_cell_58_60 ( BL60, BLN60, WL58);
sram_cell_6t_3 inst_cell_58_59 ( BL59, BLN59, WL58);
sram_cell_6t_3 inst_cell_58_58 ( BL58, BLN58, WL58);
sram_cell_6t_3 inst_cell_58_57 ( BL57, BLN57, WL58);
sram_cell_6t_3 inst_cell_58_56 ( BL56, BLN56, WL58);
sram_cell_6t_3 inst_cell_58_55 ( BL55, BLN55, WL58);
sram_cell_6t_3 inst_cell_58_54 ( BL54, BLN54, WL58);
sram_cell_6t_3 inst_cell_58_53 ( BL53, BLN53, WL58);
sram_cell_6t_3 inst_cell_58_52 ( BL52, BLN52, WL58);
sram_cell_6t_3 inst_cell_58_51 ( BL51, BLN51, WL58);
sram_cell_6t_3 inst_cell_58_50 ( BL50, BLN50, WL58);
sram_cell_6t_3 inst_cell_58_49 ( BL49, BLN49, WL58);
sram_cell_6t_3 inst_cell_58_48 ( BL48, BLN48, WL58);
sram_cell_6t_3 inst_cell_58_47 ( BL47, BLN47, WL58);
sram_cell_6t_3 inst_cell_58_46 ( BL46, BLN46, WL58);
sram_cell_6t_3 inst_cell_58_45 ( BL45, BLN45, WL58);
sram_cell_6t_3 inst_cell_58_44 ( BL44, BLN44, WL58);
sram_cell_6t_3 inst_cell_58_43 ( BL43, BLN43, WL58);
sram_cell_6t_3 inst_cell_58_42 ( BL42, BLN42, WL58);
sram_cell_6t_3 inst_cell_58_41 ( BL41, BLN41, WL58);
sram_cell_6t_3 inst_cell_58_40 ( BL40, BLN40, WL58);
sram_cell_6t_3 inst_cell_58_39 ( BL39, BLN39, WL58);
sram_cell_6t_3 inst_cell_58_38 ( BL38, BLN38, WL58);
sram_cell_6t_3 inst_cell_58_37 ( BL37, BLN37, WL58);
sram_cell_6t_3 inst_cell_58_36 ( BL36, BLN36, WL58);
sram_cell_6t_3 inst_cell_58_35 ( BL35, BLN35, WL58);
sram_cell_6t_3 inst_cell_58_34 ( BL34, BLN34, WL58);
sram_cell_6t_3 inst_cell_58_33 ( BL33, BLN33, WL58);
sram_cell_6t_3 inst_cell_58_32 ( BL32, BLN32, WL58);
sram_cell_6t_3 inst_cell_58_31 ( BL31, BLN31, WL58);
sram_cell_6t_3 inst_cell_58_30 ( BL30, BLN30, WL58);
sram_cell_6t_3 inst_cell_58_29 ( BL29, BLN29, WL58);
sram_cell_6t_3 inst_cell_58_28 ( BL28, BLN28, WL58);
sram_cell_6t_3 inst_cell_58_27 ( BL27, BLN27, WL58);
sram_cell_6t_3 inst_cell_58_26 ( BL26, BLN26, WL58);
sram_cell_6t_3 inst_cell_58_25 ( BL25, BLN25, WL58);
sram_cell_6t_3 inst_cell_58_24 ( BL24, BLN24, WL58);
sram_cell_6t_3 inst_cell_58_23 ( BL23, BLN23, WL58);
sram_cell_6t_3 inst_cell_58_22 ( BL22, BLN22, WL58);
sram_cell_6t_3 inst_cell_58_21 ( BL21, BLN21, WL58);
sram_cell_6t_3 inst_cell_58_20 ( BL20, BLN20, WL58);
sram_cell_6t_3 inst_cell_58_19 ( BL19, BLN19, WL58);
sram_cell_6t_3 inst_cell_58_18 ( BL18, BLN18, WL58);
sram_cell_6t_3 inst_cell_58_17 ( BL17, BLN17, WL58);
sram_cell_6t_3 inst_cell_58_16 ( BL16, BLN16, WL58);
sram_cell_6t_3 inst_cell_58_15 ( BL15, BLN15, WL58);
sram_cell_6t_3 inst_cell_58_14 ( BL14, BLN14, WL58);
sram_cell_6t_3 inst_cell_58_13 ( BL13, BLN13, WL58);
sram_cell_6t_3 inst_cell_58_12 ( BL12, BLN12, WL58);
sram_cell_6t_3 inst_cell_58_11 ( BL11, BLN11, WL58);
sram_cell_6t_3 inst_cell_58_10 ( BL10, BLN10, WL58);
sram_cell_6t_3 inst_cell_58_9 ( BL9, BLN9, WL58);
sram_cell_6t_3 inst_cell_58_8 ( BL8, BLN8, WL58);
sram_cell_6t_3 inst_cell_58_7 ( BL7, BLN7, WL58);
sram_cell_6t_3 inst_cell_58_6 ( BL6, BLN6, WL58);
sram_cell_6t_3 inst_cell_58_5 ( BL5, BLN5, WL58);
sram_cell_6t_3 inst_cell_58_4 ( BL4, BLN4, WL58);
sram_cell_6t_3 inst_cell_58_3 ( BL3, BLN3, WL58);
sram_cell_6t_3 inst_cell_58_2 ( BL2, BLN2, WL58);
sram_cell_6t_3 inst_cell_58_1 ( BL1, BLN1, WL58);
sram_cell_6t_3 inst_cell_58_0 ( BL0, BLN0, WL58);
sram_cell_6t_3 inst_cell_57_127 ( BL127, BLN127, WL57);
sram_cell_6t_3 inst_cell_57_126 ( BL126, BLN126, WL57);
sram_cell_6t_3 inst_cell_57_125 ( BL125, BLN125, WL57);
sram_cell_6t_3 inst_cell_57_124 ( BL124, BLN124, WL57);
sram_cell_6t_3 inst_cell_57_123 ( BL123, BLN123, WL57);
sram_cell_6t_3 inst_cell_57_122 ( BL122, BLN122, WL57);
sram_cell_6t_3 inst_cell_57_121 ( BL121, BLN121, WL57);
sram_cell_6t_3 inst_cell_57_120 ( BL120, BLN120, WL57);
sram_cell_6t_3 inst_cell_57_119 ( BL119, BLN119, WL57);
sram_cell_6t_3 inst_cell_57_118 ( BL118, BLN118, WL57);
sram_cell_6t_3 inst_cell_57_117 ( BL117, BLN117, WL57);
sram_cell_6t_3 inst_cell_57_116 ( BL116, BLN116, WL57);
sram_cell_6t_3 inst_cell_57_115 ( BL115, BLN115, WL57);
sram_cell_6t_3 inst_cell_57_114 ( BL114, BLN114, WL57);
sram_cell_6t_3 inst_cell_57_113 ( BL113, BLN113, WL57);
sram_cell_6t_3 inst_cell_57_112 ( BL112, BLN112, WL57);
sram_cell_6t_3 inst_cell_57_111 ( BL111, BLN111, WL57);
sram_cell_6t_3 inst_cell_57_110 ( BL110, BLN110, WL57);
sram_cell_6t_3 inst_cell_57_109 ( BL109, BLN109, WL57);
sram_cell_6t_3 inst_cell_57_108 ( BL108, BLN108, WL57);
sram_cell_6t_3 inst_cell_57_107 ( BL107, BLN107, WL57);
sram_cell_6t_3 inst_cell_57_106 ( BL106, BLN106, WL57);
sram_cell_6t_3 inst_cell_57_105 ( BL105, BLN105, WL57);
sram_cell_6t_3 inst_cell_57_104 ( BL104, BLN104, WL57);
sram_cell_6t_3 inst_cell_57_103 ( BL103, BLN103, WL57);
sram_cell_6t_3 inst_cell_57_102 ( BL102, BLN102, WL57);
sram_cell_6t_3 inst_cell_57_101 ( BL101, BLN101, WL57);
sram_cell_6t_3 inst_cell_57_100 ( BL100, BLN100, WL57);
sram_cell_6t_3 inst_cell_57_99 ( BL99, BLN99, WL57);
sram_cell_6t_3 inst_cell_57_98 ( BL98, BLN98, WL57);
sram_cell_6t_3 inst_cell_57_97 ( BL97, BLN97, WL57);
sram_cell_6t_3 inst_cell_57_96 ( BL96, BLN96, WL57);
sram_cell_6t_3 inst_cell_57_95 ( BL95, BLN95, WL57);
sram_cell_6t_3 inst_cell_57_94 ( BL94, BLN94, WL57);
sram_cell_6t_3 inst_cell_57_93 ( BL93, BLN93, WL57);
sram_cell_6t_3 inst_cell_57_92 ( BL92, BLN92, WL57);
sram_cell_6t_3 inst_cell_57_91 ( BL91, BLN91, WL57);
sram_cell_6t_3 inst_cell_57_90 ( BL90, BLN90, WL57);
sram_cell_6t_3 inst_cell_57_89 ( BL89, BLN89, WL57);
sram_cell_6t_3 inst_cell_57_88 ( BL88, BLN88, WL57);
sram_cell_6t_3 inst_cell_57_87 ( BL87, BLN87, WL57);
sram_cell_6t_3 inst_cell_57_86 ( BL86, BLN86, WL57);
sram_cell_6t_3 inst_cell_57_85 ( BL85, BLN85, WL57);
sram_cell_6t_3 inst_cell_57_84 ( BL84, BLN84, WL57);
sram_cell_6t_3 inst_cell_57_83 ( BL83, BLN83, WL57);
sram_cell_6t_3 inst_cell_57_82 ( BL82, BLN82, WL57);
sram_cell_6t_3 inst_cell_57_81 ( BL81, BLN81, WL57);
sram_cell_6t_3 inst_cell_57_80 ( BL80, BLN80, WL57);
sram_cell_6t_3 inst_cell_57_79 ( BL79, BLN79, WL57);
sram_cell_6t_3 inst_cell_57_78 ( BL78, BLN78, WL57);
sram_cell_6t_3 inst_cell_57_77 ( BL77, BLN77, WL57);
sram_cell_6t_3 inst_cell_57_76 ( BL76, BLN76, WL57);
sram_cell_6t_3 inst_cell_57_75 ( BL75, BLN75, WL57);
sram_cell_6t_3 inst_cell_57_74 ( BL74, BLN74, WL57);
sram_cell_6t_3 inst_cell_57_73 ( BL73, BLN73, WL57);
sram_cell_6t_3 inst_cell_57_72 ( BL72, BLN72, WL57);
sram_cell_6t_3 inst_cell_57_71 ( BL71, BLN71, WL57);
sram_cell_6t_3 inst_cell_57_70 ( BL70, BLN70, WL57);
sram_cell_6t_3 inst_cell_57_69 ( BL69, BLN69, WL57);
sram_cell_6t_3 inst_cell_57_68 ( BL68, BLN68, WL57);
sram_cell_6t_3 inst_cell_57_67 ( BL67, BLN67, WL57);
sram_cell_6t_3 inst_cell_57_66 ( BL66, BLN66, WL57);
sram_cell_6t_3 inst_cell_57_65 ( BL65, BLN65, WL57);
sram_cell_6t_3 inst_cell_57_64 ( BL64, BLN64, WL57);
sram_cell_6t_3 inst_cell_57_63 ( BL63, BLN63, WL57);
sram_cell_6t_3 inst_cell_57_62 ( BL62, BLN62, WL57);
sram_cell_6t_3 inst_cell_57_61 ( BL61, BLN61, WL57);
sram_cell_6t_3 inst_cell_57_60 ( BL60, BLN60, WL57);
sram_cell_6t_3 inst_cell_57_59 ( BL59, BLN59, WL57);
sram_cell_6t_3 inst_cell_57_58 ( BL58, BLN58, WL57);
sram_cell_6t_3 inst_cell_57_57 ( BL57, BLN57, WL57);
sram_cell_6t_3 inst_cell_57_56 ( BL56, BLN56, WL57);
sram_cell_6t_3 inst_cell_57_55 ( BL55, BLN55, WL57);
sram_cell_6t_3 inst_cell_57_54 ( BL54, BLN54, WL57);
sram_cell_6t_3 inst_cell_57_53 ( BL53, BLN53, WL57);
sram_cell_6t_3 inst_cell_57_52 ( BL52, BLN52, WL57);
sram_cell_6t_3 inst_cell_57_51 ( BL51, BLN51, WL57);
sram_cell_6t_3 inst_cell_57_50 ( BL50, BLN50, WL57);
sram_cell_6t_3 inst_cell_57_49 ( BL49, BLN49, WL57);
sram_cell_6t_3 inst_cell_57_48 ( BL48, BLN48, WL57);
sram_cell_6t_3 inst_cell_57_47 ( BL47, BLN47, WL57);
sram_cell_6t_3 inst_cell_57_46 ( BL46, BLN46, WL57);
sram_cell_6t_3 inst_cell_57_45 ( BL45, BLN45, WL57);
sram_cell_6t_3 inst_cell_57_44 ( BL44, BLN44, WL57);
sram_cell_6t_3 inst_cell_57_43 ( BL43, BLN43, WL57);
sram_cell_6t_3 inst_cell_57_42 ( BL42, BLN42, WL57);
sram_cell_6t_3 inst_cell_57_41 ( BL41, BLN41, WL57);
sram_cell_6t_3 inst_cell_57_40 ( BL40, BLN40, WL57);
sram_cell_6t_3 inst_cell_57_39 ( BL39, BLN39, WL57);
sram_cell_6t_3 inst_cell_57_38 ( BL38, BLN38, WL57);
sram_cell_6t_3 inst_cell_57_37 ( BL37, BLN37, WL57);
sram_cell_6t_3 inst_cell_57_36 ( BL36, BLN36, WL57);
sram_cell_6t_3 inst_cell_57_35 ( BL35, BLN35, WL57);
sram_cell_6t_3 inst_cell_57_34 ( BL34, BLN34, WL57);
sram_cell_6t_3 inst_cell_57_33 ( BL33, BLN33, WL57);
sram_cell_6t_3 inst_cell_57_32 ( BL32, BLN32, WL57);
sram_cell_6t_3 inst_cell_57_31 ( BL31, BLN31, WL57);
sram_cell_6t_3 inst_cell_57_30 ( BL30, BLN30, WL57);
sram_cell_6t_3 inst_cell_57_29 ( BL29, BLN29, WL57);
sram_cell_6t_3 inst_cell_57_28 ( BL28, BLN28, WL57);
sram_cell_6t_3 inst_cell_57_27 ( BL27, BLN27, WL57);
sram_cell_6t_3 inst_cell_57_26 ( BL26, BLN26, WL57);
sram_cell_6t_3 inst_cell_57_25 ( BL25, BLN25, WL57);
sram_cell_6t_3 inst_cell_57_24 ( BL24, BLN24, WL57);
sram_cell_6t_3 inst_cell_57_23 ( BL23, BLN23, WL57);
sram_cell_6t_3 inst_cell_57_22 ( BL22, BLN22, WL57);
sram_cell_6t_3 inst_cell_57_21 ( BL21, BLN21, WL57);
sram_cell_6t_3 inst_cell_57_20 ( BL20, BLN20, WL57);
sram_cell_6t_3 inst_cell_57_19 ( BL19, BLN19, WL57);
sram_cell_6t_3 inst_cell_57_18 ( BL18, BLN18, WL57);
sram_cell_6t_3 inst_cell_57_17 ( BL17, BLN17, WL57);
sram_cell_6t_3 inst_cell_57_16 ( BL16, BLN16, WL57);
sram_cell_6t_3 inst_cell_57_15 ( BL15, BLN15, WL57);
sram_cell_6t_3 inst_cell_57_14 ( BL14, BLN14, WL57);
sram_cell_6t_3 inst_cell_57_13 ( BL13, BLN13, WL57);
sram_cell_6t_3 inst_cell_57_12 ( BL12, BLN12, WL57);
sram_cell_6t_3 inst_cell_57_11 ( BL11, BLN11, WL57);
sram_cell_6t_3 inst_cell_57_10 ( BL10, BLN10, WL57);
sram_cell_6t_3 inst_cell_57_9 ( BL9, BLN9, WL57);
sram_cell_6t_3 inst_cell_57_8 ( BL8, BLN8, WL57);
sram_cell_6t_3 inst_cell_57_7 ( BL7, BLN7, WL57);
sram_cell_6t_3 inst_cell_57_6 ( BL6, BLN6, WL57);
sram_cell_6t_3 inst_cell_57_5 ( BL5, BLN5, WL57);
sram_cell_6t_3 inst_cell_57_4 ( BL4, BLN4, WL57);
sram_cell_6t_3 inst_cell_57_3 ( BL3, BLN3, WL57);
sram_cell_6t_3 inst_cell_57_2 ( BL2, BLN2, WL57);
sram_cell_6t_3 inst_cell_57_1 ( BL1, BLN1, WL57);
sram_cell_6t_3 inst_cell_57_0 ( BL0, BLN0, WL57);
sram_cell_6t_3 inst_cell_56_127 ( BL127, BLN127, WL56);
sram_cell_6t_3 inst_cell_56_126 ( BL126, BLN126, WL56);
sram_cell_6t_3 inst_cell_56_125 ( BL125, BLN125, WL56);
sram_cell_6t_3 inst_cell_56_124 ( BL124, BLN124, WL56);
sram_cell_6t_3 inst_cell_56_123 ( BL123, BLN123, WL56);
sram_cell_6t_3 inst_cell_56_122 ( BL122, BLN122, WL56);
sram_cell_6t_3 inst_cell_56_121 ( BL121, BLN121, WL56);
sram_cell_6t_3 inst_cell_56_120 ( BL120, BLN120, WL56);
sram_cell_6t_3 inst_cell_56_119 ( BL119, BLN119, WL56);
sram_cell_6t_3 inst_cell_56_118 ( BL118, BLN118, WL56);
sram_cell_6t_3 inst_cell_56_117 ( BL117, BLN117, WL56);
sram_cell_6t_3 inst_cell_56_116 ( BL116, BLN116, WL56);
sram_cell_6t_3 inst_cell_56_115 ( BL115, BLN115, WL56);
sram_cell_6t_3 inst_cell_56_114 ( BL114, BLN114, WL56);
sram_cell_6t_3 inst_cell_56_113 ( BL113, BLN113, WL56);
sram_cell_6t_3 inst_cell_56_112 ( BL112, BLN112, WL56);
sram_cell_6t_3 inst_cell_56_111 ( BL111, BLN111, WL56);
sram_cell_6t_3 inst_cell_56_110 ( BL110, BLN110, WL56);
sram_cell_6t_3 inst_cell_56_109 ( BL109, BLN109, WL56);
sram_cell_6t_3 inst_cell_56_108 ( BL108, BLN108, WL56);
sram_cell_6t_3 inst_cell_56_107 ( BL107, BLN107, WL56);
sram_cell_6t_3 inst_cell_56_106 ( BL106, BLN106, WL56);
sram_cell_6t_3 inst_cell_56_105 ( BL105, BLN105, WL56);
sram_cell_6t_3 inst_cell_56_104 ( BL104, BLN104, WL56);
sram_cell_6t_3 inst_cell_56_103 ( BL103, BLN103, WL56);
sram_cell_6t_3 inst_cell_56_102 ( BL102, BLN102, WL56);
sram_cell_6t_3 inst_cell_56_101 ( BL101, BLN101, WL56);
sram_cell_6t_3 inst_cell_56_100 ( BL100, BLN100, WL56);
sram_cell_6t_3 inst_cell_56_99 ( BL99, BLN99, WL56);
sram_cell_6t_3 inst_cell_56_98 ( BL98, BLN98, WL56);
sram_cell_6t_3 inst_cell_56_97 ( BL97, BLN97, WL56);
sram_cell_6t_3 inst_cell_56_96 ( BL96, BLN96, WL56);
sram_cell_6t_3 inst_cell_56_95 ( BL95, BLN95, WL56);
sram_cell_6t_3 inst_cell_56_94 ( BL94, BLN94, WL56);
sram_cell_6t_3 inst_cell_56_93 ( BL93, BLN93, WL56);
sram_cell_6t_3 inst_cell_56_92 ( BL92, BLN92, WL56);
sram_cell_6t_3 inst_cell_56_91 ( BL91, BLN91, WL56);
sram_cell_6t_3 inst_cell_56_90 ( BL90, BLN90, WL56);
sram_cell_6t_3 inst_cell_56_89 ( BL89, BLN89, WL56);
sram_cell_6t_3 inst_cell_56_88 ( BL88, BLN88, WL56);
sram_cell_6t_3 inst_cell_56_87 ( BL87, BLN87, WL56);
sram_cell_6t_3 inst_cell_56_86 ( BL86, BLN86, WL56);
sram_cell_6t_3 inst_cell_56_85 ( BL85, BLN85, WL56);
sram_cell_6t_3 inst_cell_56_84 ( BL84, BLN84, WL56);
sram_cell_6t_3 inst_cell_56_83 ( BL83, BLN83, WL56);
sram_cell_6t_3 inst_cell_56_82 ( BL82, BLN82, WL56);
sram_cell_6t_3 inst_cell_56_81 ( BL81, BLN81, WL56);
sram_cell_6t_3 inst_cell_56_80 ( BL80, BLN80, WL56);
sram_cell_6t_3 inst_cell_56_79 ( BL79, BLN79, WL56);
sram_cell_6t_3 inst_cell_56_78 ( BL78, BLN78, WL56);
sram_cell_6t_3 inst_cell_56_77 ( BL77, BLN77, WL56);
sram_cell_6t_3 inst_cell_56_76 ( BL76, BLN76, WL56);
sram_cell_6t_3 inst_cell_56_75 ( BL75, BLN75, WL56);
sram_cell_6t_3 inst_cell_56_74 ( BL74, BLN74, WL56);
sram_cell_6t_3 inst_cell_56_73 ( BL73, BLN73, WL56);
sram_cell_6t_3 inst_cell_56_72 ( BL72, BLN72, WL56);
sram_cell_6t_3 inst_cell_56_71 ( BL71, BLN71, WL56);
sram_cell_6t_3 inst_cell_56_70 ( BL70, BLN70, WL56);
sram_cell_6t_3 inst_cell_56_69 ( BL69, BLN69, WL56);
sram_cell_6t_3 inst_cell_56_68 ( BL68, BLN68, WL56);
sram_cell_6t_3 inst_cell_56_67 ( BL67, BLN67, WL56);
sram_cell_6t_3 inst_cell_56_66 ( BL66, BLN66, WL56);
sram_cell_6t_3 inst_cell_56_65 ( BL65, BLN65, WL56);
sram_cell_6t_3 inst_cell_56_64 ( BL64, BLN64, WL56);
sram_cell_6t_3 inst_cell_56_63 ( BL63, BLN63, WL56);
sram_cell_6t_3 inst_cell_56_62 ( BL62, BLN62, WL56);
sram_cell_6t_3 inst_cell_56_61 ( BL61, BLN61, WL56);
sram_cell_6t_3 inst_cell_56_60 ( BL60, BLN60, WL56);
sram_cell_6t_3 inst_cell_56_59 ( BL59, BLN59, WL56);
sram_cell_6t_3 inst_cell_56_58 ( BL58, BLN58, WL56);
sram_cell_6t_3 inst_cell_56_57 ( BL57, BLN57, WL56);
sram_cell_6t_3 inst_cell_56_56 ( BL56, BLN56, WL56);
sram_cell_6t_3 inst_cell_56_55 ( BL55, BLN55, WL56);
sram_cell_6t_3 inst_cell_56_54 ( BL54, BLN54, WL56);
sram_cell_6t_3 inst_cell_56_53 ( BL53, BLN53, WL56);
sram_cell_6t_3 inst_cell_56_52 ( BL52, BLN52, WL56);
sram_cell_6t_3 inst_cell_56_51 ( BL51, BLN51, WL56);
sram_cell_6t_3 inst_cell_56_50 ( BL50, BLN50, WL56);
sram_cell_6t_3 inst_cell_56_49 ( BL49, BLN49, WL56);
sram_cell_6t_3 inst_cell_56_48 ( BL48, BLN48, WL56);
sram_cell_6t_3 inst_cell_56_47 ( BL47, BLN47, WL56);
sram_cell_6t_3 inst_cell_56_46 ( BL46, BLN46, WL56);
sram_cell_6t_3 inst_cell_56_45 ( BL45, BLN45, WL56);
sram_cell_6t_3 inst_cell_56_44 ( BL44, BLN44, WL56);
sram_cell_6t_3 inst_cell_56_43 ( BL43, BLN43, WL56);
sram_cell_6t_3 inst_cell_56_42 ( BL42, BLN42, WL56);
sram_cell_6t_3 inst_cell_56_41 ( BL41, BLN41, WL56);
sram_cell_6t_3 inst_cell_56_40 ( BL40, BLN40, WL56);
sram_cell_6t_3 inst_cell_56_39 ( BL39, BLN39, WL56);
sram_cell_6t_3 inst_cell_56_38 ( BL38, BLN38, WL56);
sram_cell_6t_3 inst_cell_56_37 ( BL37, BLN37, WL56);
sram_cell_6t_3 inst_cell_56_36 ( BL36, BLN36, WL56);
sram_cell_6t_3 inst_cell_56_35 ( BL35, BLN35, WL56);
sram_cell_6t_3 inst_cell_56_34 ( BL34, BLN34, WL56);
sram_cell_6t_3 inst_cell_56_33 ( BL33, BLN33, WL56);
sram_cell_6t_3 inst_cell_56_32 ( BL32, BLN32, WL56);
sram_cell_6t_3 inst_cell_56_31 ( BL31, BLN31, WL56);
sram_cell_6t_3 inst_cell_56_30 ( BL30, BLN30, WL56);
sram_cell_6t_3 inst_cell_56_29 ( BL29, BLN29, WL56);
sram_cell_6t_3 inst_cell_56_28 ( BL28, BLN28, WL56);
sram_cell_6t_3 inst_cell_56_27 ( BL27, BLN27, WL56);
sram_cell_6t_3 inst_cell_56_26 ( BL26, BLN26, WL56);
sram_cell_6t_3 inst_cell_56_25 ( BL25, BLN25, WL56);
sram_cell_6t_3 inst_cell_56_24 ( BL24, BLN24, WL56);
sram_cell_6t_3 inst_cell_56_23 ( BL23, BLN23, WL56);
sram_cell_6t_3 inst_cell_56_22 ( BL22, BLN22, WL56);
sram_cell_6t_3 inst_cell_56_21 ( BL21, BLN21, WL56);
sram_cell_6t_3 inst_cell_56_20 ( BL20, BLN20, WL56);
sram_cell_6t_3 inst_cell_56_19 ( BL19, BLN19, WL56);
sram_cell_6t_3 inst_cell_56_18 ( BL18, BLN18, WL56);
sram_cell_6t_3 inst_cell_56_17 ( BL17, BLN17, WL56);
sram_cell_6t_3 inst_cell_56_16 ( BL16, BLN16, WL56);
sram_cell_6t_3 inst_cell_56_15 ( BL15, BLN15, WL56);
sram_cell_6t_3 inst_cell_56_14 ( BL14, BLN14, WL56);
sram_cell_6t_3 inst_cell_56_13 ( BL13, BLN13, WL56);
sram_cell_6t_3 inst_cell_56_12 ( BL12, BLN12, WL56);
sram_cell_6t_3 inst_cell_56_11 ( BL11, BLN11, WL56);
sram_cell_6t_3 inst_cell_56_10 ( BL10, BLN10, WL56);
sram_cell_6t_3 inst_cell_56_9 ( BL9, BLN9, WL56);
sram_cell_6t_3 inst_cell_56_8 ( BL8, BLN8, WL56);
sram_cell_6t_3 inst_cell_56_7 ( BL7, BLN7, WL56);
sram_cell_6t_3 inst_cell_56_6 ( BL6, BLN6, WL56);
sram_cell_6t_3 inst_cell_56_5 ( BL5, BLN5, WL56);
sram_cell_6t_3 inst_cell_56_4 ( BL4, BLN4, WL56);
sram_cell_6t_3 inst_cell_56_3 ( BL3, BLN3, WL56);
sram_cell_6t_3 inst_cell_56_2 ( BL2, BLN2, WL56);
sram_cell_6t_3 inst_cell_56_1 ( BL1, BLN1, WL56);
sram_cell_6t_3 inst_cell_56_0 ( BL0, BLN0, WL56);
sram_cell_6t_3 inst_cell_55_127 ( BL127, BLN127, WL55);
sram_cell_6t_3 inst_cell_55_126 ( BL126, BLN126, WL55);
sram_cell_6t_3 inst_cell_55_125 ( BL125, BLN125, WL55);
sram_cell_6t_3 inst_cell_55_124 ( BL124, BLN124, WL55);
sram_cell_6t_3 inst_cell_55_123 ( BL123, BLN123, WL55);
sram_cell_6t_3 inst_cell_55_122 ( BL122, BLN122, WL55);
sram_cell_6t_3 inst_cell_55_121 ( BL121, BLN121, WL55);
sram_cell_6t_3 inst_cell_55_120 ( BL120, BLN120, WL55);
sram_cell_6t_3 inst_cell_55_119 ( BL119, BLN119, WL55);
sram_cell_6t_3 inst_cell_55_118 ( BL118, BLN118, WL55);
sram_cell_6t_3 inst_cell_55_117 ( BL117, BLN117, WL55);
sram_cell_6t_3 inst_cell_55_116 ( BL116, BLN116, WL55);
sram_cell_6t_3 inst_cell_55_115 ( BL115, BLN115, WL55);
sram_cell_6t_3 inst_cell_55_114 ( BL114, BLN114, WL55);
sram_cell_6t_3 inst_cell_55_113 ( BL113, BLN113, WL55);
sram_cell_6t_3 inst_cell_55_112 ( BL112, BLN112, WL55);
sram_cell_6t_3 inst_cell_55_111 ( BL111, BLN111, WL55);
sram_cell_6t_3 inst_cell_55_110 ( BL110, BLN110, WL55);
sram_cell_6t_3 inst_cell_55_109 ( BL109, BLN109, WL55);
sram_cell_6t_3 inst_cell_55_108 ( BL108, BLN108, WL55);
sram_cell_6t_3 inst_cell_55_107 ( BL107, BLN107, WL55);
sram_cell_6t_3 inst_cell_55_106 ( BL106, BLN106, WL55);
sram_cell_6t_3 inst_cell_55_105 ( BL105, BLN105, WL55);
sram_cell_6t_3 inst_cell_55_104 ( BL104, BLN104, WL55);
sram_cell_6t_3 inst_cell_55_103 ( BL103, BLN103, WL55);
sram_cell_6t_3 inst_cell_55_102 ( BL102, BLN102, WL55);
sram_cell_6t_3 inst_cell_55_101 ( BL101, BLN101, WL55);
sram_cell_6t_3 inst_cell_55_100 ( BL100, BLN100, WL55);
sram_cell_6t_3 inst_cell_55_99 ( BL99, BLN99, WL55);
sram_cell_6t_3 inst_cell_55_98 ( BL98, BLN98, WL55);
sram_cell_6t_3 inst_cell_55_97 ( BL97, BLN97, WL55);
sram_cell_6t_3 inst_cell_55_96 ( BL96, BLN96, WL55);
sram_cell_6t_3 inst_cell_55_95 ( BL95, BLN95, WL55);
sram_cell_6t_3 inst_cell_55_94 ( BL94, BLN94, WL55);
sram_cell_6t_3 inst_cell_55_93 ( BL93, BLN93, WL55);
sram_cell_6t_3 inst_cell_55_92 ( BL92, BLN92, WL55);
sram_cell_6t_3 inst_cell_55_91 ( BL91, BLN91, WL55);
sram_cell_6t_3 inst_cell_55_90 ( BL90, BLN90, WL55);
sram_cell_6t_3 inst_cell_55_89 ( BL89, BLN89, WL55);
sram_cell_6t_3 inst_cell_55_88 ( BL88, BLN88, WL55);
sram_cell_6t_3 inst_cell_55_87 ( BL87, BLN87, WL55);
sram_cell_6t_3 inst_cell_55_86 ( BL86, BLN86, WL55);
sram_cell_6t_3 inst_cell_55_85 ( BL85, BLN85, WL55);
sram_cell_6t_3 inst_cell_55_84 ( BL84, BLN84, WL55);
sram_cell_6t_3 inst_cell_55_83 ( BL83, BLN83, WL55);
sram_cell_6t_3 inst_cell_55_82 ( BL82, BLN82, WL55);
sram_cell_6t_3 inst_cell_55_81 ( BL81, BLN81, WL55);
sram_cell_6t_3 inst_cell_55_80 ( BL80, BLN80, WL55);
sram_cell_6t_3 inst_cell_55_79 ( BL79, BLN79, WL55);
sram_cell_6t_3 inst_cell_55_78 ( BL78, BLN78, WL55);
sram_cell_6t_3 inst_cell_55_77 ( BL77, BLN77, WL55);
sram_cell_6t_3 inst_cell_55_76 ( BL76, BLN76, WL55);
sram_cell_6t_3 inst_cell_55_75 ( BL75, BLN75, WL55);
sram_cell_6t_3 inst_cell_55_74 ( BL74, BLN74, WL55);
sram_cell_6t_3 inst_cell_55_73 ( BL73, BLN73, WL55);
sram_cell_6t_3 inst_cell_55_72 ( BL72, BLN72, WL55);
sram_cell_6t_3 inst_cell_55_71 ( BL71, BLN71, WL55);
sram_cell_6t_3 inst_cell_55_70 ( BL70, BLN70, WL55);
sram_cell_6t_3 inst_cell_55_69 ( BL69, BLN69, WL55);
sram_cell_6t_3 inst_cell_55_68 ( BL68, BLN68, WL55);
sram_cell_6t_3 inst_cell_55_67 ( BL67, BLN67, WL55);
sram_cell_6t_3 inst_cell_55_66 ( BL66, BLN66, WL55);
sram_cell_6t_3 inst_cell_55_65 ( BL65, BLN65, WL55);
sram_cell_6t_3 inst_cell_55_64 ( BL64, BLN64, WL55);
sram_cell_6t_3 inst_cell_55_63 ( BL63, BLN63, WL55);
sram_cell_6t_3 inst_cell_55_62 ( BL62, BLN62, WL55);
sram_cell_6t_3 inst_cell_55_61 ( BL61, BLN61, WL55);
sram_cell_6t_3 inst_cell_55_60 ( BL60, BLN60, WL55);
sram_cell_6t_3 inst_cell_55_59 ( BL59, BLN59, WL55);
sram_cell_6t_3 inst_cell_55_58 ( BL58, BLN58, WL55);
sram_cell_6t_3 inst_cell_55_57 ( BL57, BLN57, WL55);
sram_cell_6t_3 inst_cell_55_56 ( BL56, BLN56, WL55);
sram_cell_6t_3 inst_cell_55_55 ( BL55, BLN55, WL55);
sram_cell_6t_3 inst_cell_55_54 ( BL54, BLN54, WL55);
sram_cell_6t_3 inst_cell_55_53 ( BL53, BLN53, WL55);
sram_cell_6t_3 inst_cell_55_52 ( BL52, BLN52, WL55);
sram_cell_6t_3 inst_cell_55_51 ( BL51, BLN51, WL55);
sram_cell_6t_3 inst_cell_55_50 ( BL50, BLN50, WL55);
sram_cell_6t_3 inst_cell_55_49 ( BL49, BLN49, WL55);
sram_cell_6t_3 inst_cell_55_48 ( BL48, BLN48, WL55);
sram_cell_6t_3 inst_cell_55_47 ( BL47, BLN47, WL55);
sram_cell_6t_3 inst_cell_55_46 ( BL46, BLN46, WL55);
sram_cell_6t_3 inst_cell_55_45 ( BL45, BLN45, WL55);
sram_cell_6t_3 inst_cell_55_44 ( BL44, BLN44, WL55);
sram_cell_6t_3 inst_cell_55_43 ( BL43, BLN43, WL55);
sram_cell_6t_3 inst_cell_55_42 ( BL42, BLN42, WL55);
sram_cell_6t_3 inst_cell_55_41 ( BL41, BLN41, WL55);
sram_cell_6t_3 inst_cell_55_40 ( BL40, BLN40, WL55);
sram_cell_6t_3 inst_cell_55_39 ( BL39, BLN39, WL55);
sram_cell_6t_3 inst_cell_55_38 ( BL38, BLN38, WL55);
sram_cell_6t_3 inst_cell_55_37 ( BL37, BLN37, WL55);
sram_cell_6t_3 inst_cell_55_36 ( BL36, BLN36, WL55);
sram_cell_6t_3 inst_cell_55_35 ( BL35, BLN35, WL55);
sram_cell_6t_3 inst_cell_55_34 ( BL34, BLN34, WL55);
sram_cell_6t_3 inst_cell_55_33 ( BL33, BLN33, WL55);
sram_cell_6t_3 inst_cell_55_32 ( BL32, BLN32, WL55);
sram_cell_6t_3 inst_cell_55_31 ( BL31, BLN31, WL55);
sram_cell_6t_3 inst_cell_55_30 ( BL30, BLN30, WL55);
sram_cell_6t_3 inst_cell_55_29 ( BL29, BLN29, WL55);
sram_cell_6t_3 inst_cell_55_28 ( BL28, BLN28, WL55);
sram_cell_6t_3 inst_cell_55_27 ( BL27, BLN27, WL55);
sram_cell_6t_3 inst_cell_55_26 ( BL26, BLN26, WL55);
sram_cell_6t_3 inst_cell_55_25 ( BL25, BLN25, WL55);
sram_cell_6t_3 inst_cell_55_24 ( BL24, BLN24, WL55);
sram_cell_6t_3 inst_cell_55_23 ( BL23, BLN23, WL55);
sram_cell_6t_3 inst_cell_55_22 ( BL22, BLN22, WL55);
sram_cell_6t_3 inst_cell_55_21 ( BL21, BLN21, WL55);
sram_cell_6t_3 inst_cell_55_20 ( BL20, BLN20, WL55);
sram_cell_6t_3 inst_cell_55_19 ( BL19, BLN19, WL55);
sram_cell_6t_3 inst_cell_55_18 ( BL18, BLN18, WL55);
sram_cell_6t_3 inst_cell_55_17 ( BL17, BLN17, WL55);
sram_cell_6t_3 inst_cell_55_16 ( BL16, BLN16, WL55);
sram_cell_6t_3 inst_cell_55_15 ( BL15, BLN15, WL55);
sram_cell_6t_3 inst_cell_55_14 ( BL14, BLN14, WL55);
sram_cell_6t_3 inst_cell_55_13 ( BL13, BLN13, WL55);
sram_cell_6t_3 inst_cell_55_12 ( BL12, BLN12, WL55);
sram_cell_6t_3 inst_cell_55_11 ( BL11, BLN11, WL55);
sram_cell_6t_3 inst_cell_55_10 ( BL10, BLN10, WL55);
sram_cell_6t_3 inst_cell_55_9 ( BL9, BLN9, WL55);
sram_cell_6t_3 inst_cell_55_8 ( BL8, BLN8, WL55);
sram_cell_6t_3 inst_cell_55_7 ( BL7, BLN7, WL55);
sram_cell_6t_3 inst_cell_55_6 ( BL6, BLN6, WL55);
sram_cell_6t_3 inst_cell_55_5 ( BL5, BLN5, WL55);
sram_cell_6t_3 inst_cell_55_4 ( BL4, BLN4, WL55);
sram_cell_6t_3 inst_cell_55_3 ( BL3, BLN3, WL55);
sram_cell_6t_3 inst_cell_55_2 ( BL2, BLN2, WL55);
sram_cell_6t_3 inst_cell_55_1 ( BL1, BLN1, WL55);
sram_cell_6t_3 inst_cell_55_0 ( BL0, BLN0, WL55);
sram_cell_6t_3 inst_cell_54_127 ( BL127, BLN127, WL54);
sram_cell_6t_3 inst_cell_54_126 ( BL126, BLN126, WL54);
sram_cell_6t_3 inst_cell_54_125 ( BL125, BLN125, WL54);
sram_cell_6t_3 inst_cell_54_124 ( BL124, BLN124, WL54);
sram_cell_6t_3 inst_cell_54_123 ( BL123, BLN123, WL54);
sram_cell_6t_3 inst_cell_54_122 ( BL122, BLN122, WL54);
sram_cell_6t_3 inst_cell_54_121 ( BL121, BLN121, WL54);
sram_cell_6t_3 inst_cell_54_120 ( BL120, BLN120, WL54);
sram_cell_6t_3 inst_cell_54_119 ( BL119, BLN119, WL54);
sram_cell_6t_3 inst_cell_54_118 ( BL118, BLN118, WL54);
sram_cell_6t_3 inst_cell_54_117 ( BL117, BLN117, WL54);
sram_cell_6t_3 inst_cell_54_116 ( BL116, BLN116, WL54);
sram_cell_6t_3 inst_cell_54_115 ( BL115, BLN115, WL54);
sram_cell_6t_3 inst_cell_54_114 ( BL114, BLN114, WL54);
sram_cell_6t_3 inst_cell_54_113 ( BL113, BLN113, WL54);
sram_cell_6t_3 inst_cell_54_112 ( BL112, BLN112, WL54);
sram_cell_6t_3 inst_cell_54_111 ( BL111, BLN111, WL54);
sram_cell_6t_3 inst_cell_54_110 ( BL110, BLN110, WL54);
sram_cell_6t_3 inst_cell_54_109 ( BL109, BLN109, WL54);
sram_cell_6t_3 inst_cell_54_108 ( BL108, BLN108, WL54);
sram_cell_6t_3 inst_cell_54_107 ( BL107, BLN107, WL54);
sram_cell_6t_3 inst_cell_54_106 ( BL106, BLN106, WL54);
sram_cell_6t_3 inst_cell_54_105 ( BL105, BLN105, WL54);
sram_cell_6t_3 inst_cell_54_104 ( BL104, BLN104, WL54);
sram_cell_6t_3 inst_cell_54_103 ( BL103, BLN103, WL54);
sram_cell_6t_3 inst_cell_54_102 ( BL102, BLN102, WL54);
sram_cell_6t_3 inst_cell_54_101 ( BL101, BLN101, WL54);
sram_cell_6t_3 inst_cell_54_100 ( BL100, BLN100, WL54);
sram_cell_6t_3 inst_cell_54_99 ( BL99, BLN99, WL54);
sram_cell_6t_3 inst_cell_54_98 ( BL98, BLN98, WL54);
sram_cell_6t_3 inst_cell_54_97 ( BL97, BLN97, WL54);
sram_cell_6t_3 inst_cell_54_96 ( BL96, BLN96, WL54);
sram_cell_6t_3 inst_cell_54_95 ( BL95, BLN95, WL54);
sram_cell_6t_3 inst_cell_54_94 ( BL94, BLN94, WL54);
sram_cell_6t_3 inst_cell_54_93 ( BL93, BLN93, WL54);
sram_cell_6t_3 inst_cell_54_92 ( BL92, BLN92, WL54);
sram_cell_6t_3 inst_cell_54_91 ( BL91, BLN91, WL54);
sram_cell_6t_3 inst_cell_54_90 ( BL90, BLN90, WL54);
sram_cell_6t_3 inst_cell_54_89 ( BL89, BLN89, WL54);
sram_cell_6t_3 inst_cell_54_88 ( BL88, BLN88, WL54);
sram_cell_6t_3 inst_cell_54_87 ( BL87, BLN87, WL54);
sram_cell_6t_3 inst_cell_54_86 ( BL86, BLN86, WL54);
sram_cell_6t_3 inst_cell_54_85 ( BL85, BLN85, WL54);
sram_cell_6t_3 inst_cell_54_84 ( BL84, BLN84, WL54);
sram_cell_6t_3 inst_cell_54_83 ( BL83, BLN83, WL54);
sram_cell_6t_3 inst_cell_54_82 ( BL82, BLN82, WL54);
sram_cell_6t_3 inst_cell_54_81 ( BL81, BLN81, WL54);
sram_cell_6t_3 inst_cell_54_80 ( BL80, BLN80, WL54);
sram_cell_6t_3 inst_cell_54_79 ( BL79, BLN79, WL54);
sram_cell_6t_3 inst_cell_54_78 ( BL78, BLN78, WL54);
sram_cell_6t_3 inst_cell_54_77 ( BL77, BLN77, WL54);
sram_cell_6t_3 inst_cell_54_76 ( BL76, BLN76, WL54);
sram_cell_6t_3 inst_cell_54_75 ( BL75, BLN75, WL54);
sram_cell_6t_3 inst_cell_54_74 ( BL74, BLN74, WL54);
sram_cell_6t_3 inst_cell_54_73 ( BL73, BLN73, WL54);
sram_cell_6t_3 inst_cell_54_72 ( BL72, BLN72, WL54);
sram_cell_6t_3 inst_cell_54_71 ( BL71, BLN71, WL54);
sram_cell_6t_3 inst_cell_54_70 ( BL70, BLN70, WL54);
sram_cell_6t_3 inst_cell_54_69 ( BL69, BLN69, WL54);
sram_cell_6t_3 inst_cell_54_68 ( BL68, BLN68, WL54);
sram_cell_6t_3 inst_cell_54_67 ( BL67, BLN67, WL54);
sram_cell_6t_3 inst_cell_54_66 ( BL66, BLN66, WL54);
sram_cell_6t_3 inst_cell_54_65 ( BL65, BLN65, WL54);
sram_cell_6t_3 inst_cell_54_64 ( BL64, BLN64, WL54);
sram_cell_6t_3 inst_cell_54_63 ( BL63, BLN63, WL54);
sram_cell_6t_3 inst_cell_54_62 ( BL62, BLN62, WL54);
sram_cell_6t_3 inst_cell_54_61 ( BL61, BLN61, WL54);
sram_cell_6t_3 inst_cell_54_60 ( BL60, BLN60, WL54);
sram_cell_6t_3 inst_cell_54_59 ( BL59, BLN59, WL54);
sram_cell_6t_3 inst_cell_54_58 ( BL58, BLN58, WL54);
sram_cell_6t_3 inst_cell_54_57 ( BL57, BLN57, WL54);
sram_cell_6t_3 inst_cell_54_56 ( BL56, BLN56, WL54);
sram_cell_6t_3 inst_cell_54_55 ( BL55, BLN55, WL54);
sram_cell_6t_3 inst_cell_54_54 ( BL54, BLN54, WL54);
sram_cell_6t_3 inst_cell_54_53 ( BL53, BLN53, WL54);
sram_cell_6t_3 inst_cell_54_52 ( BL52, BLN52, WL54);
sram_cell_6t_3 inst_cell_54_51 ( BL51, BLN51, WL54);
sram_cell_6t_3 inst_cell_54_50 ( BL50, BLN50, WL54);
sram_cell_6t_3 inst_cell_54_49 ( BL49, BLN49, WL54);
sram_cell_6t_3 inst_cell_54_48 ( BL48, BLN48, WL54);
sram_cell_6t_3 inst_cell_54_47 ( BL47, BLN47, WL54);
sram_cell_6t_3 inst_cell_54_46 ( BL46, BLN46, WL54);
sram_cell_6t_3 inst_cell_54_45 ( BL45, BLN45, WL54);
sram_cell_6t_3 inst_cell_54_44 ( BL44, BLN44, WL54);
sram_cell_6t_3 inst_cell_54_43 ( BL43, BLN43, WL54);
sram_cell_6t_3 inst_cell_54_42 ( BL42, BLN42, WL54);
sram_cell_6t_3 inst_cell_54_41 ( BL41, BLN41, WL54);
sram_cell_6t_3 inst_cell_54_40 ( BL40, BLN40, WL54);
sram_cell_6t_3 inst_cell_54_39 ( BL39, BLN39, WL54);
sram_cell_6t_3 inst_cell_54_38 ( BL38, BLN38, WL54);
sram_cell_6t_3 inst_cell_54_37 ( BL37, BLN37, WL54);
sram_cell_6t_3 inst_cell_54_36 ( BL36, BLN36, WL54);
sram_cell_6t_3 inst_cell_54_35 ( BL35, BLN35, WL54);
sram_cell_6t_3 inst_cell_54_34 ( BL34, BLN34, WL54);
sram_cell_6t_3 inst_cell_54_33 ( BL33, BLN33, WL54);
sram_cell_6t_3 inst_cell_54_32 ( BL32, BLN32, WL54);
sram_cell_6t_3 inst_cell_54_31 ( BL31, BLN31, WL54);
sram_cell_6t_3 inst_cell_54_30 ( BL30, BLN30, WL54);
sram_cell_6t_3 inst_cell_54_29 ( BL29, BLN29, WL54);
sram_cell_6t_3 inst_cell_54_28 ( BL28, BLN28, WL54);
sram_cell_6t_3 inst_cell_54_27 ( BL27, BLN27, WL54);
sram_cell_6t_3 inst_cell_54_26 ( BL26, BLN26, WL54);
sram_cell_6t_3 inst_cell_54_25 ( BL25, BLN25, WL54);
sram_cell_6t_3 inst_cell_54_24 ( BL24, BLN24, WL54);
sram_cell_6t_3 inst_cell_54_23 ( BL23, BLN23, WL54);
sram_cell_6t_3 inst_cell_54_22 ( BL22, BLN22, WL54);
sram_cell_6t_3 inst_cell_54_21 ( BL21, BLN21, WL54);
sram_cell_6t_3 inst_cell_54_20 ( BL20, BLN20, WL54);
sram_cell_6t_3 inst_cell_54_19 ( BL19, BLN19, WL54);
sram_cell_6t_3 inst_cell_54_18 ( BL18, BLN18, WL54);
sram_cell_6t_3 inst_cell_54_17 ( BL17, BLN17, WL54);
sram_cell_6t_3 inst_cell_54_16 ( BL16, BLN16, WL54);
sram_cell_6t_3 inst_cell_54_15 ( BL15, BLN15, WL54);
sram_cell_6t_3 inst_cell_54_14 ( BL14, BLN14, WL54);
sram_cell_6t_3 inst_cell_54_13 ( BL13, BLN13, WL54);
sram_cell_6t_3 inst_cell_54_12 ( BL12, BLN12, WL54);
sram_cell_6t_3 inst_cell_54_11 ( BL11, BLN11, WL54);
sram_cell_6t_3 inst_cell_54_10 ( BL10, BLN10, WL54);
sram_cell_6t_3 inst_cell_54_9 ( BL9, BLN9, WL54);
sram_cell_6t_3 inst_cell_54_8 ( BL8, BLN8, WL54);
sram_cell_6t_3 inst_cell_54_7 ( BL7, BLN7, WL54);
sram_cell_6t_3 inst_cell_54_6 ( BL6, BLN6, WL54);
sram_cell_6t_3 inst_cell_54_5 ( BL5, BLN5, WL54);
sram_cell_6t_3 inst_cell_54_4 ( BL4, BLN4, WL54);
sram_cell_6t_3 inst_cell_54_3 ( BL3, BLN3, WL54);
sram_cell_6t_3 inst_cell_54_2 ( BL2, BLN2, WL54);
sram_cell_6t_3 inst_cell_54_1 ( BL1, BLN1, WL54);
sram_cell_6t_3 inst_cell_54_0 ( BL0, BLN0, WL54);
sram_cell_6t_3 inst_cell_53_127 ( BL127, BLN127, WL53);
sram_cell_6t_3 inst_cell_53_126 ( BL126, BLN126, WL53);
sram_cell_6t_3 inst_cell_53_125 ( BL125, BLN125, WL53);
sram_cell_6t_3 inst_cell_53_124 ( BL124, BLN124, WL53);
sram_cell_6t_3 inst_cell_53_123 ( BL123, BLN123, WL53);
sram_cell_6t_3 inst_cell_53_122 ( BL122, BLN122, WL53);
sram_cell_6t_3 inst_cell_53_121 ( BL121, BLN121, WL53);
sram_cell_6t_3 inst_cell_53_120 ( BL120, BLN120, WL53);
sram_cell_6t_3 inst_cell_53_119 ( BL119, BLN119, WL53);
sram_cell_6t_3 inst_cell_53_118 ( BL118, BLN118, WL53);
sram_cell_6t_3 inst_cell_53_117 ( BL117, BLN117, WL53);
sram_cell_6t_3 inst_cell_53_116 ( BL116, BLN116, WL53);
sram_cell_6t_3 inst_cell_53_115 ( BL115, BLN115, WL53);
sram_cell_6t_3 inst_cell_53_114 ( BL114, BLN114, WL53);
sram_cell_6t_3 inst_cell_53_113 ( BL113, BLN113, WL53);
sram_cell_6t_3 inst_cell_53_112 ( BL112, BLN112, WL53);
sram_cell_6t_3 inst_cell_53_111 ( BL111, BLN111, WL53);
sram_cell_6t_3 inst_cell_53_110 ( BL110, BLN110, WL53);
sram_cell_6t_3 inst_cell_53_109 ( BL109, BLN109, WL53);
sram_cell_6t_3 inst_cell_53_108 ( BL108, BLN108, WL53);
sram_cell_6t_3 inst_cell_53_107 ( BL107, BLN107, WL53);
sram_cell_6t_3 inst_cell_53_106 ( BL106, BLN106, WL53);
sram_cell_6t_3 inst_cell_53_105 ( BL105, BLN105, WL53);
sram_cell_6t_3 inst_cell_53_104 ( BL104, BLN104, WL53);
sram_cell_6t_3 inst_cell_53_103 ( BL103, BLN103, WL53);
sram_cell_6t_3 inst_cell_53_102 ( BL102, BLN102, WL53);
sram_cell_6t_3 inst_cell_53_101 ( BL101, BLN101, WL53);
sram_cell_6t_3 inst_cell_53_100 ( BL100, BLN100, WL53);
sram_cell_6t_3 inst_cell_53_99 ( BL99, BLN99, WL53);
sram_cell_6t_3 inst_cell_53_98 ( BL98, BLN98, WL53);
sram_cell_6t_3 inst_cell_53_97 ( BL97, BLN97, WL53);
sram_cell_6t_3 inst_cell_53_96 ( BL96, BLN96, WL53);
sram_cell_6t_3 inst_cell_53_95 ( BL95, BLN95, WL53);
sram_cell_6t_3 inst_cell_53_94 ( BL94, BLN94, WL53);
sram_cell_6t_3 inst_cell_53_93 ( BL93, BLN93, WL53);
sram_cell_6t_3 inst_cell_53_92 ( BL92, BLN92, WL53);
sram_cell_6t_3 inst_cell_53_91 ( BL91, BLN91, WL53);
sram_cell_6t_3 inst_cell_53_90 ( BL90, BLN90, WL53);
sram_cell_6t_3 inst_cell_53_89 ( BL89, BLN89, WL53);
sram_cell_6t_3 inst_cell_53_88 ( BL88, BLN88, WL53);
sram_cell_6t_3 inst_cell_53_87 ( BL87, BLN87, WL53);
sram_cell_6t_3 inst_cell_53_86 ( BL86, BLN86, WL53);
sram_cell_6t_3 inst_cell_53_85 ( BL85, BLN85, WL53);
sram_cell_6t_3 inst_cell_53_84 ( BL84, BLN84, WL53);
sram_cell_6t_3 inst_cell_53_83 ( BL83, BLN83, WL53);
sram_cell_6t_3 inst_cell_53_82 ( BL82, BLN82, WL53);
sram_cell_6t_3 inst_cell_53_81 ( BL81, BLN81, WL53);
sram_cell_6t_3 inst_cell_53_80 ( BL80, BLN80, WL53);
sram_cell_6t_3 inst_cell_53_79 ( BL79, BLN79, WL53);
sram_cell_6t_3 inst_cell_53_78 ( BL78, BLN78, WL53);
sram_cell_6t_3 inst_cell_53_77 ( BL77, BLN77, WL53);
sram_cell_6t_3 inst_cell_53_76 ( BL76, BLN76, WL53);
sram_cell_6t_3 inst_cell_53_75 ( BL75, BLN75, WL53);
sram_cell_6t_3 inst_cell_53_74 ( BL74, BLN74, WL53);
sram_cell_6t_3 inst_cell_53_73 ( BL73, BLN73, WL53);
sram_cell_6t_3 inst_cell_53_72 ( BL72, BLN72, WL53);
sram_cell_6t_3 inst_cell_53_71 ( BL71, BLN71, WL53);
sram_cell_6t_3 inst_cell_53_70 ( BL70, BLN70, WL53);
sram_cell_6t_3 inst_cell_53_69 ( BL69, BLN69, WL53);
sram_cell_6t_3 inst_cell_53_68 ( BL68, BLN68, WL53);
sram_cell_6t_3 inst_cell_53_67 ( BL67, BLN67, WL53);
sram_cell_6t_3 inst_cell_53_66 ( BL66, BLN66, WL53);
sram_cell_6t_3 inst_cell_53_65 ( BL65, BLN65, WL53);
sram_cell_6t_3 inst_cell_53_64 ( BL64, BLN64, WL53);
sram_cell_6t_3 inst_cell_53_63 ( BL63, BLN63, WL53);
sram_cell_6t_3 inst_cell_53_62 ( BL62, BLN62, WL53);
sram_cell_6t_3 inst_cell_53_61 ( BL61, BLN61, WL53);
sram_cell_6t_3 inst_cell_53_60 ( BL60, BLN60, WL53);
sram_cell_6t_3 inst_cell_53_59 ( BL59, BLN59, WL53);
sram_cell_6t_3 inst_cell_53_58 ( BL58, BLN58, WL53);
sram_cell_6t_3 inst_cell_53_57 ( BL57, BLN57, WL53);
sram_cell_6t_3 inst_cell_53_56 ( BL56, BLN56, WL53);
sram_cell_6t_3 inst_cell_53_55 ( BL55, BLN55, WL53);
sram_cell_6t_3 inst_cell_53_54 ( BL54, BLN54, WL53);
sram_cell_6t_3 inst_cell_53_53 ( BL53, BLN53, WL53);
sram_cell_6t_3 inst_cell_53_52 ( BL52, BLN52, WL53);
sram_cell_6t_3 inst_cell_53_51 ( BL51, BLN51, WL53);
sram_cell_6t_3 inst_cell_53_50 ( BL50, BLN50, WL53);
sram_cell_6t_3 inst_cell_53_49 ( BL49, BLN49, WL53);
sram_cell_6t_3 inst_cell_53_48 ( BL48, BLN48, WL53);
sram_cell_6t_3 inst_cell_53_47 ( BL47, BLN47, WL53);
sram_cell_6t_3 inst_cell_53_46 ( BL46, BLN46, WL53);
sram_cell_6t_3 inst_cell_53_45 ( BL45, BLN45, WL53);
sram_cell_6t_3 inst_cell_53_44 ( BL44, BLN44, WL53);
sram_cell_6t_3 inst_cell_53_43 ( BL43, BLN43, WL53);
sram_cell_6t_3 inst_cell_53_42 ( BL42, BLN42, WL53);
sram_cell_6t_3 inst_cell_53_41 ( BL41, BLN41, WL53);
sram_cell_6t_3 inst_cell_53_40 ( BL40, BLN40, WL53);
sram_cell_6t_3 inst_cell_53_39 ( BL39, BLN39, WL53);
sram_cell_6t_3 inst_cell_53_38 ( BL38, BLN38, WL53);
sram_cell_6t_3 inst_cell_53_37 ( BL37, BLN37, WL53);
sram_cell_6t_3 inst_cell_53_36 ( BL36, BLN36, WL53);
sram_cell_6t_3 inst_cell_53_35 ( BL35, BLN35, WL53);
sram_cell_6t_3 inst_cell_53_34 ( BL34, BLN34, WL53);
sram_cell_6t_3 inst_cell_53_33 ( BL33, BLN33, WL53);
sram_cell_6t_3 inst_cell_53_32 ( BL32, BLN32, WL53);
sram_cell_6t_3 inst_cell_53_31 ( BL31, BLN31, WL53);
sram_cell_6t_3 inst_cell_53_30 ( BL30, BLN30, WL53);
sram_cell_6t_3 inst_cell_53_29 ( BL29, BLN29, WL53);
sram_cell_6t_3 inst_cell_53_28 ( BL28, BLN28, WL53);
sram_cell_6t_3 inst_cell_53_27 ( BL27, BLN27, WL53);
sram_cell_6t_3 inst_cell_53_26 ( BL26, BLN26, WL53);
sram_cell_6t_3 inst_cell_53_25 ( BL25, BLN25, WL53);
sram_cell_6t_3 inst_cell_53_24 ( BL24, BLN24, WL53);
sram_cell_6t_3 inst_cell_53_23 ( BL23, BLN23, WL53);
sram_cell_6t_3 inst_cell_53_22 ( BL22, BLN22, WL53);
sram_cell_6t_3 inst_cell_53_21 ( BL21, BLN21, WL53);
sram_cell_6t_3 inst_cell_53_20 ( BL20, BLN20, WL53);
sram_cell_6t_3 inst_cell_53_19 ( BL19, BLN19, WL53);
sram_cell_6t_3 inst_cell_53_18 ( BL18, BLN18, WL53);
sram_cell_6t_3 inst_cell_53_17 ( BL17, BLN17, WL53);
sram_cell_6t_3 inst_cell_53_16 ( BL16, BLN16, WL53);
sram_cell_6t_3 inst_cell_53_15 ( BL15, BLN15, WL53);
sram_cell_6t_3 inst_cell_53_14 ( BL14, BLN14, WL53);
sram_cell_6t_3 inst_cell_53_13 ( BL13, BLN13, WL53);
sram_cell_6t_3 inst_cell_53_12 ( BL12, BLN12, WL53);
sram_cell_6t_3 inst_cell_53_11 ( BL11, BLN11, WL53);
sram_cell_6t_3 inst_cell_53_10 ( BL10, BLN10, WL53);
sram_cell_6t_3 inst_cell_53_9 ( BL9, BLN9, WL53);
sram_cell_6t_3 inst_cell_53_8 ( BL8, BLN8, WL53);
sram_cell_6t_3 inst_cell_53_7 ( BL7, BLN7, WL53);
sram_cell_6t_3 inst_cell_53_6 ( BL6, BLN6, WL53);
sram_cell_6t_3 inst_cell_53_5 ( BL5, BLN5, WL53);
sram_cell_6t_3 inst_cell_53_4 ( BL4, BLN4, WL53);
sram_cell_6t_3 inst_cell_53_3 ( BL3, BLN3, WL53);
sram_cell_6t_3 inst_cell_53_2 ( BL2, BLN2, WL53);
sram_cell_6t_3 inst_cell_53_1 ( BL1, BLN1, WL53);
sram_cell_6t_3 inst_cell_53_0 ( BL0, BLN0, WL53);
sram_cell_6t_3 inst_cell_52_127 ( BL127, BLN127, WL52);
sram_cell_6t_3 inst_cell_52_126 ( BL126, BLN126, WL52);
sram_cell_6t_3 inst_cell_52_125 ( BL125, BLN125, WL52);
sram_cell_6t_3 inst_cell_52_124 ( BL124, BLN124, WL52);
sram_cell_6t_3 inst_cell_52_123 ( BL123, BLN123, WL52);
sram_cell_6t_3 inst_cell_52_122 ( BL122, BLN122, WL52);
sram_cell_6t_3 inst_cell_52_121 ( BL121, BLN121, WL52);
sram_cell_6t_3 inst_cell_52_120 ( BL120, BLN120, WL52);
sram_cell_6t_3 inst_cell_52_119 ( BL119, BLN119, WL52);
sram_cell_6t_3 inst_cell_52_118 ( BL118, BLN118, WL52);
sram_cell_6t_3 inst_cell_52_117 ( BL117, BLN117, WL52);
sram_cell_6t_3 inst_cell_52_116 ( BL116, BLN116, WL52);
sram_cell_6t_3 inst_cell_52_115 ( BL115, BLN115, WL52);
sram_cell_6t_3 inst_cell_52_114 ( BL114, BLN114, WL52);
sram_cell_6t_3 inst_cell_52_113 ( BL113, BLN113, WL52);
sram_cell_6t_3 inst_cell_52_112 ( BL112, BLN112, WL52);
sram_cell_6t_3 inst_cell_52_111 ( BL111, BLN111, WL52);
sram_cell_6t_3 inst_cell_52_110 ( BL110, BLN110, WL52);
sram_cell_6t_3 inst_cell_52_109 ( BL109, BLN109, WL52);
sram_cell_6t_3 inst_cell_52_108 ( BL108, BLN108, WL52);
sram_cell_6t_3 inst_cell_52_107 ( BL107, BLN107, WL52);
sram_cell_6t_3 inst_cell_52_106 ( BL106, BLN106, WL52);
sram_cell_6t_3 inst_cell_52_105 ( BL105, BLN105, WL52);
sram_cell_6t_3 inst_cell_52_104 ( BL104, BLN104, WL52);
sram_cell_6t_3 inst_cell_52_103 ( BL103, BLN103, WL52);
sram_cell_6t_3 inst_cell_52_102 ( BL102, BLN102, WL52);
sram_cell_6t_3 inst_cell_52_101 ( BL101, BLN101, WL52);
sram_cell_6t_3 inst_cell_52_100 ( BL100, BLN100, WL52);
sram_cell_6t_3 inst_cell_52_99 ( BL99, BLN99, WL52);
sram_cell_6t_3 inst_cell_52_98 ( BL98, BLN98, WL52);
sram_cell_6t_3 inst_cell_52_97 ( BL97, BLN97, WL52);
sram_cell_6t_3 inst_cell_52_96 ( BL96, BLN96, WL52);
sram_cell_6t_3 inst_cell_52_95 ( BL95, BLN95, WL52);
sram_cell_6t_3 inst_cell_52_94 ( BL94, BLN94, WL52);
sram_cell_6t_3 inst_cell_52_93 ( BL93, BLN93, WL52);
sram_cell_6t_3 inst_cell_52_92 ( BL92, BLN92, WL52);
sram_cell_6t_3 inst_cell_52_91 ( BL91, BLN91, WL52);
sram_cell_6t_3 inst_cell_52_90 ( BL90, BLN90, WL52);
sram_cell_6t_3 inst_cell_52_89 ( BL89, BLN89, WL52);
sram_cell_6t_3 inst_cell_52_88 ( BL88, BLN88, WL52);
sram_cell_6t_3 inst_cell_52_87 ( BL87, BLN87, WL52);
sram_cell_6t_3 inst_cell_52_86 ( BL86, BLN86, WL52);
sram_cell_6t_3 inst_cell_52_85 ( BL85, BLN85, WL52);
sram_cell_6t_3 inst_cell_52_84 ( BL84, BLN84, WL52);
sram_cell_6t_3 inst_cell_52_83 ( BL83, BLN83, WL52);
sram_cell_6t_3 inst_cell_52_82 ( BL82, BLN82, WL52);
sram_cell_6t_3 inst_cell_52_81 ( BL81, BLN81, WL52);
sram_cell_6t_3 inst_cell_52_80 ( BL80, BLN80, WL52);
sram_cell_6t_3 inst_cell_52_79 ( BL79, BLN79, WL52);
sram_cell_6t_3 inst_cell_52_78 ( BL78, BLN78, WL52);
sram_cell_6t_3 inst_cell_52_77 ( BL77, BLN77, WL52);
sram_cell_6t_3 inst_cell_52_76 ( BL76, BLN76, WL52);
sram_cell_6t_3 inst_cell_52_75 ( BL75, BLN75, WL52);
sram_cell_6t_3 inst_cell_52_74 ( BL74, BLN74, WL52);
sram_cell_6t_3 inst_cell_52_73 ( BL73, BLN73, WL52);
sram_cell_6t_3 inst_cell_52_72 ( BL72, BLN72, WL52);
sram_cell_6t_3 inst_cell_52_71 ( BL71, BLN71, WL52);
sram_cell_6t_3 inst_cell_52_70 ( BL70, BLN70, WL52);
sram_cell_6t_3 inst_cell_52_69 ( BL69, BLN69, WL52);
sram_cell_6t_3 inst_cell_52_68 ( BL68, BLN68, WL52);
sram_cell_6t_3 inst_cell_52_67 ( BL67, BLN67, WL52);
sram_cell_6t_3 inst_cell_52_66 ( BL66, BLN66, WL52);
sram_cell_6t_3 inst_cell_52_65 ( BL65, BLN65, WL52);
sram_cell_6t_3 inst_cell_52_64 ( BL64, BLN64, WL52);
sram_cell_6t_3 inst_cell_52_63 ( BL63, BLN63, WL52);
sram_cell_6t_3 inst_cell_52_62 ( BL62, BLN62, WL52);
sram_cell_6t_3 inst_cell_52_61 ( BL61, BLN61, WL52);
sram_cell_6t_3 inst_cell_52_60 ( BL60, BLN60, WL52);
sram_cell_6t_3 inst_cell_52_59 ( BL59, BLN59, WL52);
sram_cell_6t_3 inst_cell_52_58 ( BL58, BLN58, WL52);
sram_cell_6t_3 inst_cell_52_57 ( BL57, BLN57, WL52);
sram_cell_6t_3 inst_cell_52_56 ( BL56, BLN56, WL52);
sram_cell_6t_3 inst_cell_52_55 ( BL55, BLN55, WL52);
sram_cell_6t_3 inst_cell_52_54 ( BL54, BLN54, WL52);
sram_cell_6t_3 inst_cell_52_53 ( BL53, BLN53, WL52);
sram_cell_6t_3 inst_cell_52_52 ( BL52, BLN52, WL52);
sram_cell_6t_3 inst_cell_52_51 ( BL51, BLN51, WL52);
sram_cell_6t_3 inst_cell_52_50 ( BL50, BLN50, WL52);
sram_cell_6t_3 inst_cell_52_49 ( BL49, BLN49, WL52);
sram_cell_6t_3 inst_cell_52_48 ( BL48, BLN48, WL52);
sram_cell_6t_3 inst_cell_52_47 ( BL47, BLN47, WL52);
sram_cell_6t_3 inst_cell_52_46 ( BL46, BLN46, WL52);
sram_cell_6t_3 inst_cell_52_45 ( BL45, BLN45, WL52);
sram_cell_6t_3 inst_cell_52_44 ( BL44, BLN44, WL52);
sram_cell_6t_3 inst_cell_52_43 ( BL43, BLN43, WL52);
sram_cell_6t_3 inst_cell_52_42 ( BL42, BLN42, WL52);
sram_cell_6t_3 inst_cell_52_41 ( BL41, BLN41, WL52);
sram_cell_6t_3 inst_cell_52_40 ( BL40, BLN40, WL52);
sram_cell_6t_3 inst_cell_52_39 ( BL39, BLN39, WL52);
sram_cell_6t_3 inst_cell_52_38 ( BL38, BLN38, WL52);
sram_cell_6t_3 inst_cell_52_37 ( BL37, BLN37, WL52);
sram_cell_6t_3 inst_cell_52_36 ( BL36, BLN36, WL52);
sram_cell_6t_3 inst_cell_52_35 ( BL35, BLN35, WL52);
sram_cell_6t_3 inst_cell_52_34 ( BL34, BLN34, WL52);
sram_cell_6t_3 inst_cell_52_33 ( BL33, BLN33, WL52);
sram_cell_6t_3 inst_cell_52_32 ( BL32, BLN32, WL52);
sram_cell_6t_3 inst_cell_52_31 ( BL31, BLN31, WL52);
sram_cell_6t_3 inst_cell_52_30 ( BL30, BLN30, WL52);
sram_cell_6t_3 inst_cell_52_29 ( BL29, BLN29, WL52);
sram_cell_6t_3 inst_cell_52_28 ( BL28, BLN28, WL52);
sram_cell_6t_3 inst_cell_52_27 ( BL27, BLN27, WL52);
sram_cell_6t_3 inst_cell_52_26 ( BL26, BLN26, WL52);
sram_cell_6t_3 inst_cell_52_25 ( BL25, BLN25, WL52);
sram_cell_6t_3 inst_cell_52_24 ( BL24, BLN24, WL52);
sram_cell_6t_3 inst_cell_52_23 ( BL23, BLN23, WL52);
sram_cell_6t_3 inst_cell_52_22 ( BL22, BLN22, WL52);
sram_cell_6t_3 inst_cell_52_21 ( BL21, BLN21, WL52);
sram_cell_6t_3 inst_cell_52_20 ( BL20, BLN20, WL52);
sram_cell_6t_3 inst_cell_52_19 ( BL19, BLN19, WL52);
sram_cell_6t_3 inst_cell_52_18 ( BL18, BLN18, WL52);
sram_cell_6t_3 inst_cell_52_17 ( BL17, BLN17, WL52);
sram_cell_6t_3 inst_cell_52_16 ( BL16, BLN16, WL52);
sram_cell_6t_3 inst_cell_52_15 ( BL15, BLN15, WL52);
sram_cell_6t_3 inst_cell_52_14 ( BL14, BLN14, WL52);
sram_cell_6t_3 inst_cell_52_13 ( BL13, BLN13, WL52);
sram_cell_6t_3 inst_cell_52_12 ( BL12, BLN12, WL52);
sram_cell_6t_3 inst_cell_52_11 ( BL11, BLN11, WL52);
sram_cell_6t_3 inst_cell_52_10 ( BL10, BLN10, WL52);
sram_cell_6t_3 inst_cell_52_9 ( BL9, BLN9, WL52);
sram_cell_6t_3 inst_cell_52_8 ( BL8, BLN8, WL52);
sram_cell_6t_3 inst_cell_52_7 ( BL7, BLN7, WL52);
sram_cell_6t_3 inst_cell_52_6 ( BL6, BLN6, WL52);
sram_cell_6t_3 inst_cell_52_5 ( BL5, BLN5, WL52);
sram_cell_6t_3 inst_cell_52_4 ( BL4, BLN4, WL52);
sram_cell_6t_3 inst_cell_52_3 ( BL3, BLN3, WL52);
sram_cell_6t_3 inst_cell_52_2 ( BL2, BLN2, WL52);
sram_cell_6t_3 inst_cell_52_1 ( BL1, BLN1, WL52);
sram_cell_6t_3 inst_cell_52_0 ( BL0, BLN0, WL52);
sram_cell_6t_3 inst_cell_51_127 ( BL127, BLN127, WL51);
sram_cell_6t_3 inst_cell_51_126 ( BL126, BLN126, WL51);
sram_cell_6t_3 inst_cell_51_125 ( BL125, BLN125, WL51);
sram_cell_6t_3 inst_cell_51_124 ( BL124, BLN124, WL51);
sram_cell_6t_3 inst_cell_51_123 ( BL123, BLN123, WL51);
sram_cell_6t_3 inst_cell_51_122 ( BL122, BLN122, WL51);
sram_cell_6t_3 inst_cell_51_121 ( BL121, BLN121, WL51);
sram_cell_6t_3 inst_cell_51_120 ( BL120, BLN120, WL51);
sram_cell_6t_3 inst_cell_51_119 ( BL119, BLN119, WL51);
sram_cell_6t_3 inst_cell_51_118 ( BL118, BLN118, WL51);
sram_cell_6t_3 inst_cell_51_117 ( BL117, BLN117, WL51);
sram_cell_6t_3 inst_cell_51_116 ( BL116, BLN116, WL51);
sram_cell_6t_3 inst_cell_51_115 ( BL115, BLN115, WL51);
sram_cell_6t_3 inst_cell_51_114 ( BL114, BLN114, WL51);
sram_cell_6t_3 inst_cell_51_113 ( BL113, BLN113, WL51);
sram_cell_6t_3 inst_cell_51_112 ( BL112, BLN112, WL51);
sram_cell_6t_3 inst_cell_51_111 ( BL111, BLN111, WL51);
sram_cell_6t_3 inst_cell_51_110 ( BL110, BLN110, WL51);
sram_cell_6t_3 inst_cell_51_109 ( BL109, BLN109, WL51);
sram_cell_6t_3 inst_cell_51_108 ( BL108, BLN108, WL51);
sram_cell_6t_3 inst_cell_51_107 ( BL107, BLN107, WL51);
sram_cell_6t_3 inst_cell_51_106 ( BL106, BLN106, WL51);
sram_cell_6t_3 inst_cell_51_105 ( BL105, BLN105, WL51);
sram_cell_6t_3 inst_cell_51_104 ( BL104, BLN104, WL51);
sram_cell_6t_3 inst_cell_51_103 ( BL103, BLN103, WL51);
sram_cell_6t_3 inst_cell_51_102 ( BL102, BLN102, WL51);
sram_cell_6t_3 inst_cell_51_101 ( BL101, BLN101, WL51);
sram_cell_6t_3 inst_cell_51_100 ( BL100, BLN100, WL51);
sram_cell_6t_3 inst_cell_51_99 ( BL99, BLN99, WL51);
sram_cell_6t_3 inst_cell_51_98 ( BL98, BLN98, WL51);
sram_cell_6t_3 inst_cell_51_97 ( BL97, BLN97, WL51);
sram_cell_6t_3 inst_cell_51_96 ( BL96, BLN96, WL51);
sram_cell_6t_3 inst_cell_51_95 ( BL95, BLN95, WL51);
sram_cell_6t_3 inst_cell_51_94 ( BL94, BLN94, WL51);
sram_cell_6t_3 inst_cell_51_93 ( BL93, BLN93, WL51);
sram_cell_6t_3 inst_cell_51_92 ( BL92, BLN92, WL51);
sram_cell_6t_3 inst_cell_51_91 ( BL91, BLN91, WL51);
sram_cell_6t_3 inst_cell_51_90 ( BL90, BLN90, WL51);
sram_cell_6t_3 inst_cell_51_89 ( BL89, BLN89, WL51);
sram_cell_6t_3 inst_cell_51_88 ( BL88, BLN88, WL51);
sram_cell_6t_3 inst_cell_51_87 ( BL87, BLN87, WL51);
sram_cell_6t_3 inst_cell_51_86 ( BL86, BLN86, WL51);
sram_cell_6t_3 inst_cell_51_85 ( BL85, BLN85, WL51);
sram_cell_6t_3 inst_cell_51_84 ( BL84, BLN84, WL51);
sram_cell_6t_3 inst_cell_51_83 ( BL83, BLN83, WL51);
sram_cell_6t_3 inst_cell_51_82 ( BL82, BLN82, WL51);
sram_cell_6t_3 inst_cell_51_81 ( BL81, BLN81, WL51);
sram_cell_6t_3 inst_cell_51_80 ( BL80, BLN80, WL51);
sram_cell_6t_3 inst_cell_51_79 ( BL79, BLN79, WL51);
sram_cell_6t_3 inst_cell_51_78 ( BL78, BLN78, WL51);
sram_cell_6t_3 inst_cell_51_77 ( BL77, BLN77, WL51);
sram_cell_6t_3 inst_cell_51_76 ( BL76, BLN76, WL51);
sram_cell_6t_3 inst_cell_51_75 ( BL75, BLN75, WL51);
sram_cell_6t_3 inst_cell_51_74 ( BL74, BLN74, WL51);
sram_cell_6t_3 inst_cell_51_73 ( BL73, BLN73, WL51);
sram_cell_6t_3 inst_cell_51_72 ( BL72, BLN72, WL51);
sram_cell_6t_3 inst_cell_51_71 ( BL71, BLN71, WL51);
sram_cell_6t_3 inst_cell_51_70 ( BL70, BLN70, WL51);
sram_cell_6t_3 inst_cell_51_69 ( BL69, BLN69, WL51);
sram_cell_6t_3 inst_cell_51_68 ( BL68, BLN68, WL51);
sram_cell_6t_3 inst_cell_51_67 ( BL67, BLN67, WL51);
sram_cell_6t_3 inst_cell_51_66 ( BL66, BLN66, WL51);
sram_cell_6t_3 inst_cell_51_65 ( BL65, BLN65, WL51);
sram_cell_6t_3 inst_cell_51_64 ( BL64, BLN64, WL51);
sram_cell_6t_3 inst_cell_51_63 ( BL63, BLN63, WL51);
sram_cell_6t_3 inst_cell_51_62 ( BL62, BLN62, WL51);
sram_cell_6t_3 inst_cell_51_61 ( BL61, BLN61, WL51);
sram_cell_6t_3 inst_cell_51_60 ( BL60, BLN60, WL51);
sram_cell_6t_3 inst_cell_51_59 ( BL59, BLN59, WL51);
sram_cell_6t_3 inst_cell_51_58 ( BL58, BLN58, WL51);
sram_cell_6t_3 inst_cell_51_57 ( BL57, BLN57, WL51);
sram_cell_6t_3 inst_cell_51_56 ( BL56, BLN56, WL51);
sram_cell_6t_3 inst_cell_51_55 ( BL55, BLN55, WL51);
sram_cell_6t_3 inst_cell_51_54 ( BL54, BLN54, WL51);
sram_cell_6t_3 inst_cell_51_53 ( BL53, BLN53, WL51);
sram_cell_6t_3 inst_cell_51_52 ( BL52, BLN52, WL51);
sram_cell_6t_3 inst_cell_51_51 ( BL51, BLN51, WL51);
sram_cell_6t_3 inst_cell_51_50 ( BL50, BLN50, WL51);
sram_cell_6t_3 inst_cell_51_49 ( BL49, BLN49, WL51);
sram_cell_6t_3 inst_cell_51_48 ( BL48, BLN48, WL51);
sram_cell_6t_3 inst_cell_51_47 ( BL47, BLN47, WL51);
sram_cell_6t_3 inst_cell_51_46 ( BL46, BLN46, WL51);
sram_cell_6t_3 inst_cell_51_45 ( BL45, BLN45, WL51);
sram_cell_6t_3 inst_cell_51_44 ( BL44, BLN44, WL51);
sram_cell_6t_3 inst_cell_51_43 ( BL43, BLN43, WL51);
sram_cell_6t_3 inst_cell_51_42 ( BL42, BLN42, WL51);
sram_cell_6t_3 inst_cell_51_41 ( BL41, BLN41, WL51);
sram_cell_6t_3 inst_cell_51_40 ( BL40, BLN40, WL51);
sram_cell_6t_3 inst_cell_51_39 ( BL39, BLN39, WL51);
sram_cell_6t_3 inst_cell_51_38 ( BL38, BLN38, WL51);
sram_cell_6t_3 inst_cell_51_37 ( BL37, BLN37, WL51);
sram_cell_6t_3 inst_cell_51_36 ( BL36, BLN36, WL51);
sram_cell_6t_3 inst_cell_51_35 ( BL35, BLN35, WL51);
sram_cell_6t_3 inst_cell_51_34 ( BL34, BLN34, WL51);
sram_cell_6t_3 inst_cell_51_33 ( BL33, BLN33, WL51);
sram_cell_6t_3 inst_cell_51_32 ( BL32, BLN32, WL51);
sram_cell_6t_3 inst_cell_51_31 ( BL31, BLN31, WL51);
sram_cell_6t_3 inst_cell_51_30 ( BL30, BLN30, WL51);
sram_cell_6t_3 inst_cell_51_29 ( BL29, BLN29, WL51);
sram_cell_6t_3 inst_cell_51_28 ( BL28, BLN28, WL51);
sram_cell_6t_3 inst_cell_51_27 ( BL27, BLN27, WL51);
sram_cell_6t_3 inst_cell_51_26 ( BL26, BLN26, WL51);
sram_cell_6t_3 inst_cell_51_25 ( BL25, BLN25, WL51);
sram_cell_6t_3 inst_cell_51_24 ( BL24, BLN24, WL51);
sram_cell_6t_3 inst_cell_51_23 ( BL23, BLN23, WL51);
sram_cell_6t_3 inst_cell_51_22 ( BL22, BLN22, WL51);
sram_cell_6t_3 inst_cell_51_21 ( BL21, BLN21, WL51);
sram_cell_6t_3 inst_cell_51_20 ( BL20, BLN20, WL51);
sram_cell_6t_3 inst_cell_51_19 ( BL19, BLN19, WL51);
sram_cell_6t_3 inst_cell_51_18 ( BL18, BLN18, WL51);
sram_cell_6t_3 inst_cell_51_17 ( BL17, BLN17, WL51);
sram_cell_6t_3 inst_cell_51_16 ( BL16, BLN16, WL51);
sram_cell_6t_3 inst_cell_51_15 ( BL15, BLN15, WL51);
sram_cell_6t_3 inst_cell_51_14 ( BL14, BLN14, WL51);
sram_cell_6t_3 inst_cell_51_13 ( BL13, BLN13, WL51);
sram_cell_6t_3 inst_cell_51_12 ( BL12, BLN12, WL51);
sram_cell_6t_3 inst_cell_51_11 ( BL11, BLN11, WL51);
sram_cell_6t_3 inst_cell_51_10 ( BL10, BLN10, WL51);
sram_cell_6t_3 inst_cell_51_9 ( BL9, BLN9, WL51);
sram_cell_6t_3 inst_cell_51_8 ( BL8, BLN8, WL51);
sram_cell_6t_3 inst_cell_51_7 ( BL7, BLN7, WL51);
sram_cell_6t_3 inst_cell_51_6 ( BL6, BLN6, WL51);
sram_cell_6t_3 inst_cell_51_5 ( BL5, BLN5, WL51);
sram_cell_6t_3 inst_cell_51_4 ( BL4, BLN4, WL51);
sram_cell_6t_3 inst_cell_51_3 ( BL3, BLN3, WL51);
sram_cell_6t_3 inst_cell_51_2 ( BL2, BLN2, WL51);
sram_cell_6t_3 inst_cell_51_1 ( BL1, BLN1, WL51);
sram_cell_6t_3 inst_cell_51_0 ( BL0, BLN0, WL51);
sram_cell_6t_3 inst_cell_50_127 ( BL127, BLN127, WL50);
sram_cell_6t_3 inst_cell_50_126 ( BL126, BLN126, WL50);
sram_cell_6t_3 inst_cell_50_125 ( BL125, BLN125, WL50);
sram_cell_6t_3 inst_cell_50_124 ( BL124, BLN124, WL50);
sram_cell_6t_3 inst_cell_50_123 ( BL123, BLN123, WL50);
sram_cell_6t_3 inst_cell_50_122 ( BL122, BLN122, WL50);
sram_cell_6t_3 inst_cell_50_121 ( BL121, BLN121, WL50);
sram_cell_6t_3 inst_cell_50_120 ( BL120, BLN120, WL50);
sram_cell_6t_3 inst_cell_50_119 ( BL119, BLN119, WL50);
sram_cell_6t_3 inst_cell_50_118 ( BL118, BLN118, WL50);
sram_cell_6t_3 inst_cell_50_117 ( BL117, BLN117, WL50);
sram_cell_6t_3 inst_cell_50_116 ( BL116, BLN116, WL50);
sram_cell_6t_3 inst_cell_50_115 ( BL115, BLN115, WL50);
sram_cell_6t_3 inst_cell_50_114 ( BL114, BLN114, WL50);
sram_cell_6t_3 inst_cell_50_113 ( BL113, BLN113, WL50);
sram_cell_6t_3 inst_cell_50_112 ( BL112, BLN112, WL50);
sram_cell_6t_3 inst_cell_50_111 ( BL111, BLN111, WL50);
sram_cell_6t_3 inst_cell_50_110 ( BL110, BLN110, WL50);
sram_cell_6t_3 inst_cell_50_109 ( BL109, BLN109, WL50);
sram_cell_6t_3 inst_cell_50_108 ( BL108, BLN108, WL50);
sram_cell_6t_3 inst_cell_50_107 ( BL107, BLN107, WL50);
sram_cell_6t_3 inst_cell_50_106 ( BL106, BLN106, WL50);
sram_cell_6t_3 inst_cell_50_105 ( BL105, BLN105, WL50);
sram_cell_6t_3 inst_cell_50_104 ( BL104, BLN104, WL50);
sram_cell_6t_3 inst_cell_50_103 ( BL103, BLN103, WL50);
sram_cell_6t_3 inst_cell_50_102 ( BL102, BLN102, WL50);
sram_cell_6t_3 inst_cell_50_101 ( BL101, BLN101, WL50);
sram_cell_6t_3 inst_cell_50_100 ( BL100, BLN100, WL50);
sram_cell_6t_3 inst_cell_50_99 ( BL99, BLN99, WL50);
sram_cell_6t_3 inst_cell_50_98 ( BL98, BLN98, WL50);
sram_cell_6t_3 inst_cell_50_97 ( BL97, BLN97, WL50);
sram_cell_6t_3 inst_cell_50_96 ( BL96, BLN96, WL50);
sram_cell_6t_3 inst_cell_50_95 ( BL95, BLN95, WL50);
sram_cell_6t_3 inst_cell_50_94 ( BL94, BLN94, WL50);
sram_cell_6t_3 inst_cell_50_93 ( BL93, BLN93, WL50);
sram_cell_6t_3 inst_cell_50_92 ( BL92, BLN92, WL50);
sram_cell_6t_3 inst_cell_50_91 ( BL91, BLN91, WL50);
sram_cell_6t_3 inst_cell_50_90 ( BL90, BLN90, WL50);
sram_cell_6t_3 inst_cell_50_89 ( BL89, BLN89, WL50);
sram_cell_6t_3 inst_cell_50_88 ( BL88, BLN88, WL50);
sram_cell_6t_3 inst_cell_50_87 ( BL87, BLN87, WL50);
sram_cell_6t_3 inst_cell_50_86 ( BL86, BLN86, WL50);
sram_cell_6t_3 inst_cell_50_85 ( BL85, BLN85, WL50);
sram_cell_6t_3 inst_cell_50_84 ( BL84, BLN84, WL50);
sram_cell_6t_3 inst_cell_50_83 ( BL83, BLN83, WL50);
sram_cell_6t_3 inst_cell_50_82 ( BL82, BLN82, WL50);
sram_cell_6t_3 inst_cell_50_81 ( BL81, BLN81, WL50);
sram_cell_6t_3 inst_cell_50_80 ( BL80, BLN80, WL50);
sram_cell_6t_3 inst_cell_50_79 ( BL79, BLN79, WL50);
sram_cell_6t_3 inst_cell_50_78 ( BL78, BLN78, WL50);
sram_cell_6t_3 inst_cell_50_77 ( BL77, BLN77, WL50);
sram_cell_6t_3 inst_cell_50_76 ( BL76, BLN76, WL50);
sram_cell_6t_3 inst_cell_50_75 ( BL75, BLN75, WL50);
sram_cell_6t_3 inst_cell_50_74 ( BL74, BLN74, WL50);
sram_cell_6t_3 inst_cell_50_73 ( BL73, BLN73, WL50);
sram_cell_6t_3 inst_cell_50_72 ( BL72, BLN72, WL50);
sram_cell_6t_3 inst_cell_50_71 ( BL71, BLN71, WL50);
sram_cell_6t_3 inst_cell_50_70 ( BL70, BLN70, WL50);
sram_cell_6t_3 inst_cell_50_69 ( BL69, BLN69, WL50);
sram_cell_6t_3 inst_cell_50_68 ( BL68, BLN68, WL50);
sram_cell_6t_3 inst_cell_50_67 ( BL67, BLN67, WL50);
sram_cell_6t_3 inst_cell_50_66 ( BL66, BLN66, WL50);
sram_cell_6t_3 inst_cell_50_65 ( BL65, BLN65, WL50);
sram_cell_6t_3 inst_cell_50_64 ( BL64, BLN64, WL50);
sram_cell_6t_3 inst_cell_50_63 ( BL63, BLN63, WL50);
sram_cell_6t_3 inst_cell_50_62 ( BL62, BLN62, WL50);
sram_cell_6t_3 inst_cell_50_61 ( BL61, BLN61, WL50);
sram_cell_6t_3 inst_cell_50_60 ( BL60, BLN60, WL50);
sram_cell_6t_3 inst_cell_50_59 ( BL59, BLN59, WL50);
sram_cell_6t_3 inst_cell_50_58 ( BL58, BLN58, WL50);
sram_cell_6t_3 inst_cell_50_57 ( BL57, BLN57, WL50);
sram_cell_6t_3 inst_cell_50_56 ( BL56, BLN56, WL50);
sram_cell_6t_3 inst_cell_50_55 ( BL55, BLN55, WL50);
sram_cell_6t_3 inst_cell_50_54 ( BL54, BLN54, WL50);
sram_cell_6t_3 inst_cell_50_53 ( BL53, BLN53, WL50);
sram_cell_6t_3 inst_cell_50_52 ( BL52, BLN52, WL50);
sram_cell_6t_3 inst_cell_50_51 ( BL51, BLN51, WL50);
sram_cell_6t_3 inst_cell_50_50 ( BL50, BLN50, WL50);
sram_cell_6t_3 inst_cell_50_49 ( BL49, BLN49, WL50);
sram_cell_6t_3 inst_cell_50_48 ( BL48, BLN48, WL50);
sram_cell_6t_3 inst_cell_50_47 ( BL47, BLN47, WL50);
sram_cell_6t_3 inst_cell_50_46 ( BL46, BLN46, WL50);
sram_cell_6t_3 inst_cell_50_45 ( BL45, BLN45, WL50);
sram_cell_6t_3 inst_cell_50_44 ( BL44, BLN44, WL50);
sram_cell_6t_3 inst_cell_50_43 ( BL43, BLN43, WL50);
sram_cell_6t_3 inst_cell_50_42 ( BL42, BLN42, WL50);
sram_cell_6t_3 inst_cell_50_41 ( BL41, BLN41, WL50);
sram_cell_6t_3 inst_cell_50_40 ( BL40, BLN40, WL50);
sram_cell_6t_3 inst_cell_50_39 ( BL39, BLN39, WL50);
sram_cell_6t_3 inst_cell_50_38 ( BL38, BLN38, WL50);
sram_cell_6t_3 inst_cell_50_37 ( BL37, BLN37, WL50);
sram_cell_6t_3 inst_cell_50_36 ( BL36, BLN36, WL50);
sram_cell_6t_3 inst_cell_50_35 ( BL35, BLN35, WL50);
sram_cell_6t_3 inst_cell_50_34 ( BL34, BLN34, WL50);
sram_cell_6t_3 inst_cell_50_33 ( BL33, BLN33, WL50);
sram_cell_6t_3 inst_cell_50_32 ( BL32, BLN32, WL50);
sram_cell_6t_3 inst_cell_50_31 ( BL31, BLN31, WL50);
sram_cell_6t_3 inst_cell_50_30 ( BL30, BLN30, WL50);
sram_cell_6t_3 inst_cell_50_29 ( BL29, BLN29, WL50);
sram_cell_6t_3 inst_cell_50_28 ( BL28, BLN28, WL50);
sram_cell_6t_3 inst_cell_50_27 ( BL27, BLN27, WL50);
sram_cell_6t_3 inst_cell_50_26 ( BL26, BLN26, WL50);
sram_cell_6t_3 inst_cell_50_25 ( BL25, BLN25, WL50);
sram_cell_6t_3 inst_cell_50_24 ( BL24, BLN24, WL50);
sram_cell_6t_3 inst_cell_50_23 ( BL23, BLN23, WL50);
sram_cell_6t_3 inst_cell_50_22 ( BL22, BLN22, WL50);
sram_cell_6t_3 inst_cell_50_21 ( BL21, BLN21, WL50);
sram_cell_6t_3 inst_cell_50_20 ( BL20, BLN20, WL50);
sram_cell_6t_3 inst_cell_50_19 ( BL19, BLN19, WL50);
sram_cell_6t_3 inst_cell_50_18 ( BL18, BLN18, WL50);
sram_cell_6t_3 inst_cell_50_17 ( BL17, BLN17, WL50);
sram_cell_6t_3 inst_cell_50_16 ( BL16, BLN16, WL50);
sram_cell_6t_3 inst_cell_50_15 ( BL15, BLN15, WL50);
sram_cell_6t_3 inst_cell_50_14 ( BL14, BLN14, WL50);
sram_cell_6t_3 inst_cell_50_13 ( BL13, BLN13, WL50);
sram_cell_6t_3 inst_cell_50_12 ( BL12, BLN12, WL50);
sram_cell_6t_3 inst_cell_50_11 ( BL11, BLN11, WL50);
sram_cell_6t_3 inst_cell_50_10 ( BL10, BLN10, WL50);
sram_cell_6t_3 inst_cell_50_9 ( BL9, BLN9, WL50);
sram_cell_6t_3 inst_cell_50_8 ( BL8, BLN8, WL50);
sram_cell_6t_3 inst_cell_50_7 ( BL7, BLN7, WL50);
sram_cell_6t_3 inst_cell_50_6 ( BL6, BLN6, WL50);
sram_cell_6t_3 inst_cell_50_5 ( BL5, BLN5, WL50);
sram_cell_6t_3 inst_cell_50_4 ( BL4, BLN4, WL50);
sram_cell_6t_3 inst_cell_50_3 ( BL3, BLN3, WL50);
sram_cell_6t_3 inst_cell_50_2 ( BL2, BLN2, WL50);
sram_cell_6t_3 inst_cell_50_1 ( BL1, BLN1, WL50);
sram_cell_6t_3 inst_cell_50_0 ( BL0, BLN0, WL50);
sram_cell_6t_3 inst_cell_49_127 ( BL127, BLN127, WL49);
sram_cell_6t_3 inst_cell_49_126 ( BL126, BLN126, WL49);
sram_cell_6t_3 inst_cell_49_125 ( BL125, BLN125, WL49);
sram_cell_6t_3 inst_cell_49_124 ( BL124, BLN124, WL49);
sram_cell_6t_3 inst_cell_49_123 ( BL123, BLN123, WL49);
sram_cell_6t_3 inst_cell_49_122 ( BL122, BLN122, WL49);
sram_cell_6t_3 inst_cell_49_121 ( BL121, BLN121, WL49);
sram_cell_6t_3 inst_cell_49_120 ( BL120, BLN120, WL49);
sram_cell_6t_3 inst_cell_49_119 ( BL119, BLN119, WL49);
sram_cell_6t_3 inst_cell_49_118 ( BL118, BLN118, WL49);
sram_cell_6t_3 inst_cell_49_117 ( BL117, BLN117, WL49);
sram_cell_6t_3 inst_cell_49_116 ( BL116, BLN116, WL49);
sram_cell_6t_3 inst_cell_49_115 ( BL115, BLN115, WL49);
sram_cell_6t_3 inst_cell_49_114 ( BL114, BLN114, WL49);
sram_cell_6t_3 inst_cell_49_113 ( BL113, BLN113, WL49);
sram_cell_6t_3 inst_cell_49_112 ( BL112, BLN112, WL49);
sram_cell_6t_3 inst_cell_49_111 ( BL111, BLN111, WL49);
sram_cell_6t_3 inst_cell_49_110 ( BL110, BLN110, WL49);
sram_cell_6t_3 inst_cell_49_109 ( BL109, BLN109, WL49);
sram_cell_6t_3 inst_cell_49_108 ( BL108, BLN108, WL49);
sram_cell_6t_3 inst_cell_49_107 ( BL107, BLN107, WL49);
sram_cell_6t_3 inst_cell_49_106 ( BL106, BLN106, WL49);
sram_cell_6t_3 inst_cell_49_105 ( BL105, BLN105, WL49);
sram_cell_6t_3 inst_cell_49_104 ( BL104, BLN104, WL49);
sram_cell_6t_3 inst_cell_49_103 ( BL103, BLN103, WL49);
sram_cell_6t_3 inst_cell_49_102 ( BL102, BLN102, WL49);
sram_cell_6t_3 inst_cell_49_101 ( BL101, BLN101, WL49);
sram_cell_6t_3 inst_cell_49_100 ( BL100, BLN100, WL49);
sram_cell_6t_3 inst_cell_49_99 ( BL99, BLN99, WL49);
sram_cell_6t_3 inst_cell_49_98 ( BL98, BLN98, WL49);
sram_cell_6t_3 inst_cell_49_97 ( BL97, BLN97, WL49);
sram_cell_6t_3 inst_cell_49_96 ( BL96, BLN96, WL49);
sram_cell_6t_3 inst_cell_49_95 ( BL95, BLN95, WL49);
sram_cell_6t_3 inst_cell_49_94 ( BL94, BLN94, WL49);
sram_cell_6t_3 inst_cell_49_93 ( BL93, BLN93, WL49);
sram_cell_6t_3 inst_cell_49_92 ( BL92, BLN92, WL49);
sram_cell_6t_3 inst_cell_49_91 ( BL91, BLN91, WL49);
sram_cell_6t_3 inst_cell_49_90 ( BL90, BLN90, WL49);
sram_cell_6t_3 inst_cell_49_89 ( BL89, BLN89, WL49);
sram_cell_6t_3 inst_cell_49_88 ( BL88, BLN88, WL49);
sram_cell_6t_3 inst_cell_49_87 ( BL87, BLN87, WL49);
sram_cell_6t_3 inst_cell_49_86 ( BL86, BLN86, WL49);
sram_cell_6t_3 inst_cell_49_85 ( BL85, BLN85, WL49);
sram_cell_6t_3 inst_cell_49_84 ( BL84, BLN84, WL49);
sram_cell_6t_3 inst_cell_49_83 ( BL83, BLN83, WL49);
sram_cell_6t_3 inst_cell_49_82 ( BL82, BLN82, WL49);
sram_cell_6t_3 inst_cell_49_81 ( BL81, BLN81, WL49);
sram_cell_6t_3 inst_cell_49_80 ( BL80, BLN80, WL49);
sram_cell_6t_3 inst_cell_49_79 ( BL79, BLN79, WL49);
sram_cell_6t_3 inst_cell_49_78 ( BL78, BLN78, WL49);
sram_cell_6t_3 inst_cell_49_77 ( BL77, BLN77, WL49);
sram_cell_6t_3 inst_cell_49_76 ( BL76, BLN76, WL49);
sram_cell_6t_3 inst_cell_49_75 ( BL75, BLN75, WL49);
sram_cell_6t_3 inst_cell_49_74 ( BL74, BLN74, WL49);
sram_cell_6t_3 inst_cell_49_73 ( BL73, BLN73, WL49);
sram_cell_6t_3 inst_cell_49_72 ( BL72, BLN72, WL49);
sram_cell_6t_3 inst_cell_49_71 ( BL71, BLN71, WL49);
sram_cell_6t_3 inst_cell_49_70 ( BL70, BLN70, WL49);
sram_cell_6t_3 inst_cell_49_69 ( BL69, BLN69, WL49);
sram_cell_6t_3 inst_cell_49_68 ( BL68, BLN68, WL49);
sram_cell_6t_3 inst_cell_49_67 ( BL67, BLN67, WL49);
sram_cell_6t_3 inst_cell_49_66 ( BL66, BLN66, WL49);
sram_cell_6t_3 inst_cell_49_65 ( BL65, BLN65, WL49);
sram_cell_6t_3 inst_cell_49_64 ( BL64, BLN64, WL49);
sram_cell_6t_3 inst_cell_49_63 ( BL63, BLN63, WL49);
sram_cell_6t_3 inst_cell_49_62 ( BL62, BLN62, WL49);
sram_cell_6t_3 inst_cell_49_61 ( BL61, BLN61, WL49);
sram_cell_6t_3 inst_cell_49_60 ( BL60, BLN60, WL49);
sram_cell_6t_3 inst_cell_49_59 ( BL59, BLN59, WL49);
sram_cell_6t_3 inst_cell_49_58 ( BL58, BLN58, WL49);
sram_cell_6t_3 inst_cell_49_57 ( BL57, BLN57, WL49);
sram_cell_6t_3 inst_cell_49_56 ( BL56, BLN56, WL49);
sram_cell_6t_3 inst_cell_49_55 ( BL55, BLN55, WL49);
sram_cell_6t_3 inst_cell_49_54 ( BL54, BLN54, WL49);
sram_cell_6t_3 inst_cell_49_53 ( BL53, BLN53, WL49);
sram_cell_6t_3 inst_cell_49_52 ( BL52, BLN52, WL49);
sram_cell_6t_3 inst_cell_49_51 ( BL51, BLN51, WL49);
sram_cell_6t_3 inst_cell_49_50 ( BL50, BLN50, WL49);
sram_cell_6t_3 inst_cell_49_49 ( BL49, BLN49, WL49);
sram_cell_6t_3 inst_cell_49_48 ( BL48, BLN48, WL49);
sram_cell_6t_3 inst_cell_49_47 ( BL47, BLN47, WL49);
sram_cell_6t_3 inst_cell_49_46 ( BL46, BLN46, WL49);
sram_cell_6t_3 inst_cell_49_45 ( BL45, BLN45, WL49);
sram_cell_6t_3 inst_cell_49_44 ( BL44, BLN44, WL49);
sram_cell_6t_3 inst_cell_49_43 ( BL43, BLN43, WL49);
sram_cell_6t_3 inst_cell_49_42 ( BL42, BLN42, WL49);
sram_cell_6t_3 inst_cell_49_41 ( BL41, BLN41, WL49);
sram_cell_6t_3 inst_cell_49_40 ( BL40, BLN40, WL49);
sram_cell_6t_3 inst_cell_49_39 ( BL39, BLN39, WL49);
sram_cell_6t_3 inst_cell_49_38 ( BL38, BLN38, WL49);
sram_cell_6t_3 inst_cell_49_37 ( BL37, BLN37, WL49);
sram_cell_6t_3 inst_cell_49_36 ( BL36, BLN36, WL49);
sram_cell_6t_3 inst_cell_49_35 ( BL35, BLN35, WL49);
sram_cell_6t_3 inst_cell_49_34 ( BL34, BLN34, WL49);
sram_cell_6t_3 inst_cell_49_33 ( BL33, BLN33, WL49);
sram_cell_6t_3 inst_cell_49_32 ( BL32, BLN32, WL49);
sram_cell_6t_3 inst_cell_49_31 ( BL31, BLN31, WL49);
sram_cell_6t_3 inst_cell_49_30 ( BL30, BLN30, WL49);
sram_cell_6t_3 inst_cell_49_29 ( BL29, BLN29, WL49);
sram_cell_6t_3 inst_cell_49_28 ( BL28, BLN28, WL49);
sram_cell_6t_3 inst_cell_49_27 ( BL27, BLN27, WL49);
sram_cell_6t_3 inst_cell_49_26 ( BL26, BLN26, WL49);
sram_cell_6t_3 inst_cell_49_25 ( BL25, BLN25, WL49);
sram_cell_6t_3 inst_cell_49_24 ( BL24, BLN24, WL49);
sram_cell_6t_3 inst_cell_49_23 ( BL23, BLN23, WL49);
sram_cell_6t_3 inst_cell_49_22 ( BL22, BLN22, WL49);
sram_cell_6t_3 inst_cell_49_21 ( BL21, BLN21, WL49);
sram_cell_6t_3 inst_cell_49_20 ( BL20, BLN20, WL49);
sram_cell_6t_3 inst_cell_49_19 ( BL19, BLN19, WL49);
sram_cell_6t_3 inst_cell_49_18 ( BL18, BLN18, WL49);
sram_cell_6t_3 inst_cell_49_17 ( BL17, BLN17, WL49);
sram_cell_6t_3 inst_cell_49_16 ( BL16, BLN16, WL49);
sram_cell_6t_3 inst_cell_49_15 ( BL15, BLN15, WL49);
sram_cell_6t_3 inst_cell_49_14 ( BL14, BLN14, WL49);
sram_cell_6t_3 inst_cell_49_13 ( BL13, BLN13, WL49);
sram_cell_6t_3 inst_cell_49_12 ( BL12, BLN12, WL49);
sram_cell_6t_3 inst_cell_49_11 ( BL11, BLN11, WL49);
sram_cell_6t_3 inst_cell_49_10 ( BL10, BLN10, WL49);
sram_cell_6t_3 inst_cell_49_9 ( BL9, BLN9, WL49);
sram_cell_6t_3 inst_cell_49_8 ( BL8, BLN8, WL49);
sram_cell_6t_3 inst_cell_49_7 ( BL7, BLN7, WL49);
sram_cell_6t_3 inst_cell_49_6 ( BL6, BLN6, WL49);
sram_cell_6t_3 inst_cell_49_5 ( BL5, BLN5, WL49);
sram_cell_6t_3 inst_cell_49_4 ( BL4, BLN4, WL49);
sram_cell_6t_3 inst_cell_49_3 ( BL3, BLN3, WL49);
sram_cell_6t_3 inst_cell_49_2 ( BL2, BLN2, WL49);
sram_cell_6t_3 inst_cell_49_1 ( BL1, BLN1, WL49);
sram_cell_6t_3 inst_cell_49_0 ( BL0, BLN0, WL49);
sram_cell_6t_3 inst_cell_48_127 ( BL127, BLN127, WL48);
sram_cell_6t_3 inst_cell_48_126 ( BL126, BLN126, WL48);
sram_cell_6t_3 inst_cell_48_125 ( BL125, BLN125, WL48);
sram_cell_6t_3 inst_cell_48_124 ( BL124, BLN124, WL48);
sram_cell_6t_3 inst_cell_48_123 ( BL123, BLN123, WL48);
sram_cell_6t_3 inst_cell_48_122 ( BL122, BLN122, WL48);
sram_cell_6t_3 inst_cell_48_121 ( BL121, BLN121, WL48);
sram_cell_6t_3 inst_cell_48_120 ( BL120, BLN120, WL48);
sram_cell_6t_3 inst_cell_48_119 ( BL119, BLN119, WL48);
sram_cell_6t_3 inst_cell_48_118 ( BL118, BLN118, WL48);
sram_cell_6t_3 inst_cell_48_117 ( BL117, BLN117, WL48);
sram_cell_6t_3 inst_cell_48_116 ( BL116, BLN116, WL48);
sram_cell_6t_3 inst_cell_48_115 ( BL115, BLN115, WL48);
sram_cell_6t_3 inst_cell_48_114 ( BL114, BLN114, WL48);
sram_cell_6t_3 inst_cell_48_113 ( BL113, BLN113, WL48);
sram_cell_6t_3 inst_cell_48_112 ( BL112, BLN112, WL48);
sram_cell_6t_3 inst_cell_48_111 ( BL111, BLN111, WL48);
sram_cell_6t_3 inst_cell_48_110 ( BL110, BLN110, WL48);
sram_cell_6t_3 inst_cell_48_109 ( BL109, BLN109, WL48);
sram_cell_6t_3 inst_cell_48_108 ( BL108, BLN108, WL48);
sram_cell_6t_3 inst_cell_48_107 ( BL107, BLN107, WL48);
sram_cell_6t_3 inst_cell_48_106 ( BL106, BLN106, WL48);
sram_cell_6t_3 inst_cell_48_105 ( BL105, BLN105, WL48);
sram_cell_6t_3 inst_cell_48_104 ( BL104, BLN104, WL48);
sram_cell_6t_3 inst_cell_48_103 ( BL103, BLN103, WL48);
sram_cell_6t_3 inst_cell_48_102 ( BL102, BLN102, WL48);
sram_cell_6t_3 inst_cell_48_101 ( BL101, BLN101, WL48);
sram_cell_6t_3 inst_cell_48_100 ( BL100, BLN100, WL48);
sram_cell_6t_3 inst_cell_48_99 ( BL99, BLN99, WL48);
sram_cell_6t_3 inst_cell_48_98 ( BL98, BLN98, WL48);
sram_cell_6t_3 inst_cell_48_97 ( BL97, BLN97, WL48);
sram_cell_6t_3 inst_cell_48_96 ( BL96, BLN96, WL48);
sram_cell_6t_3 inst_cell_48_95 ( BL95, BLN95, WL48);
sram_cell_6t_3 inst_cell_48_94 ( BL94, BLN94, WL48);
sram_cell_6t_3 inst_cell_48_93 ( BL93, BLN93, WL48);
sram_cell_6t_3 inst_cell_48_92 ( BL92, BLN92, WL48);
sram_cell_6t_3 inst_cell_48_91 ( BL91, BLN91, WL48);
sram_cell_6t_3 inst_cell_48_90 ( BL90, BLN90, WL48);
sram_cell_6t_3 inst_cell_48_89 ( BL89, BLN89, WL48);
sram_cell_6t_3 inst_cell_48_88 ( BL88, BLN88, WL48);
sram_cell_6t_3 inst_cell_48_87 ( BL87, BLN87, WL48);
sram_cell_6t_3 inst_cell_48_86 ( BL86, BLN86, WL48);
sram_cell_6t_3 inst_cell_48_85 ( BL85, BLN85, WL48);
sram_cell_6t_3 inst_cell_48_84 ( BL84, BLN84, WL48);
sram_cell_6t_3 inst_cell_48_83 ( BL83, BLN83, WL48);
sram_cell_6t_3 inst_cell_48_82 ( BL82, BLN82, WL48);
sram_cell_6t_3 inst_cell_48_81 ( BL81, BLN81, WL48);
sram_cell_6t_3 inst_cell_48_80 ( BL80, BLN80, WL48);
sram_cell_6t_3 inst_cell_48_79 ( BL79, BLN79, WL48);
sram_cell_6t_3 inst_cell_48_78 ( BL78, BLN78, WL48);
sram_cell_6t_3 inst_cell_48_77 ( BL77, BLN77, WL48);
sram_cell_6t_3 inst_cell_48_76 ( BL76, BLN76, WL48);
sram_cell_6t_3 inst_cell_48_75 ( BL75, BLN75, WL48);
sram_cell_6t_3 inst_cell_48_74 ( BL74, BLN74, WL48);
sram_cell_6t_3 inst_cell_48_73 ( BL73, BLN73, WL48);
sram_cell_6t_3 inst_cell_48_72 ( BL72, BLN72, WL48);
sram_cell_6t_3 inst_cell_48_71 ( BL71, BLN71, WL48);
sram_cell_6t_3 inst_cell_48_70 ( BL70, BLN70, WL48);
sram_cell_6t_3 inst_cell_48_69 ( BL69, BLN69, WL48);
sram_cell_6t_3 inst_cell_48_68 ( BL68, BLN68, WL48);
sram_cell_6t_3 inst_cell_48_67 ( BL67, BLN67, WL48);
sram_cell_6t_3 inst_cell_48_66 ( BL66, BLN66, WL48);
sram_cell_6t_3 inst_cell_48_65 ( BL65, BLN65, WL48);
sram_cell_6t_3 inst_cell_48_64 ( BL64, BLN64, WL48);
sram_cell_6t_3 inst_cell_48_63 ( BL63, BLN63, WL48);
sram_cell_6t_3 inst_cell_48_62 ( BL62, BLN62, WL48);
sram_cell_6t_3 inst_cell_48_61 ( BL61, BLN61, WL48);
sram_cell_6t_3 inst_cell_48_60 ( BL60, BLN60, WL48);
sram_cell_6t_3 inst_cell_48_59 ( BL59, BLN59, WL48);
sram_cell_6t_3 inst_cell_48_58 ( BL58, BLN58, WL48);
sram_cell_6t_3 inst_cell_48_57 ( BL57, BLN57, WL48);
sram_cell_6t_3 inst_cell_48_56 ( BL56, BLN56, WL48);
sram_cell_6t_3 inst_cell_48_55 ( BL55, BLN55, WL48);
sram_cell_6t_3 inst_cell_48_54 ( BL54, BLN54, WL48);
sram_cell_6t_3 inst_cell_48_53 ( BL53, BLN53, WL48);
sram_cell_6t_3 inst_cell_48_52 ( BL52, BLN52, WL48);
sram_cell_6t_3 inst_cell_48_51 ( BL51, BLN51, WL48);
sram_cell_6t_3 inst_cell_48_50 ( BL50, BLN50, WL48);
sram_cell_6t_3 inst_cell_48_49 ( BL49, BLN49, WL48);
sram_cell_6t_3 inst_cell_48_48 ( BL48, BLN48, WL48);
sram_cell_6t_3 inst_cell_48_47 ( BL47, BLN47, WL48);
sram_cell_6t_3 inst_cell_48_46 ( BL46, BLN46, WL48);
sram_cell_6t_3 inst_cell_48_45 ( BL45, BLN45, WL48);
sram_cell_6t_3 inst_cell_48_44 ( BL44, BLN44, WL48);
sram_cell_6t_3 inst_cell_48_43 ( BL43, BLN43, WL48);
sram_cell_6t_3 inst_cell_48_42 ( BL42, BLN42, WL48);
sram_cell_6t_3 inst_cell_48_41 ( BL41, BLN41, WL48);
sram_cell_6t_3 inst_cell_48_40 ( BL40, BLN40, WL48);
sram_cell_6t_3 inst_cell_48_39 ( BL39, BLN39, WL48);
sram_cell_6t_3 inst_cell_48_38 ( BL38, BLN38, WL48);
sram_cell_6t_3 inst_cell_48_37 ( BL37, BLN37, WL48);
sram_cell_6t_3 inst_cell_48_36 ( BL36, BLN36, WL48);
sram_cell_6t_3 inst_cell_48_35 ( BL35, BLN35, WL48);
sram_cell_6t_3 inst_cell_48_34 ( BL34, BLN34, WL48);
sram_cell_6t_3 inst_cell_48_33 ( BL33, BLN33, WL48);
sram_cell_6t_3 inst_cell_48_32 ( BL32, BLN32, WL48);
sram_cell_6t_3 inst_cell_48_31 ( BL31, BLN31, WL48);
sram_cell_6t_3 inst_cell_48_30 ( BL30, BLN30, WL48);
sram_cell_6t_3 inst_cell_48_29 ( BL29, BLN29, WL48);
sram_cell_6t_3 inst_cell_48_28 ( BL28, BLN28, WL48);
sram_cell_6t_3 inst_cell_48_27 ( BL27, BLN27, WL48);
sram_cell_6t_3 inst_cell_48_26 ( BL26, BLN26, WL48);
sram_cell_6t_3 inst_cell_48_25 ( BL25, BLN25, WL48);
sram_cell_6t_3 inst_cell_48_24 ( BL24, BLN24, WL48);
sram_cell_6t_3 inst_cell_48_23 ( BL23, BLN23, WL48);
sram_cell_6t_3 inst_cell_48_22 ( BL22, BLN22, WL48);
sram_cell_6t_3 inst_cell_48_21 ( BL21, BLN21, WL48);
sram_cell_6t_3 inst_cell_48_20 ( BL20, BLN20, WL48);
sram_cell_6t_3 inst_cell_48_19 ( BL19, BLN19, WL48);
sram_cell_6t_3 inst_cell_48_18 ( BL18, BLN18, WL48);
sram_cell_6t_3 inst_cell_48_17 ( BL17, BLN17, WL48);
sram_cell_6t_3 inst_cell_48_16 ( BL16, BLN16, WL48);
sram_cell_6t_3 inst_cell_48_15 ( BL15, BLN15, WL48);
sram_cell_6t_3 inst_cell_48_14 ( BL14, BLN14, WL48);
sram_cell_6t_3 inst_cell_48_13 ( BL13, BLN13, WL48);
sram_cell_6t_3 inst_cell_48_12 ( BL12, BLN12, WL48);
sram_cell_6t_3 inst_cell_48_11 ( BL11, BLN11, WL48);
sram_cell_6t_3 inst_cell_48_10 ( BL10, BLN10, WL48);
sram_cell_6t_3 inst_cell_48_9 ( BL9, BLN9, WL48);
sram_cell_6t_3 inst_cell_48_8 ( BL8, BLN8, WL48);
sram_cell_6t_3 inst_cell_48_7 ( BL7, BLN7, WL48);
sram_cell_6t_3 inst_cell_48_6 ( BL6, BLN6, WL48);
sram_cell_6t_3 inst_cell_48_5 ( BL5, BLN5, WL48);
sram_cell_6t_3 inst_cell_48_4 ( BL4, BLN4, WL48);
sram_cell_6t_3 inst_cell_48_3 ( BL3, BLN3, WL48);
sram_cell_6t_3 inst_cell_48_2 ( BL2, BLN2, WL48);
sram_cell_6t_3 inst_cell_48_1 ( BL1, BLN1, WL48);
sram_cell_6t_3 inst_cell_48_0 ( BL0, BLN0, WL48);
sram_cell_6t_3 inst_cell_47_127 ( BL127, BLN127, WL47);
sram_cell_6t_3 inst_cell_47_126 ( BL126, BLN126, WL47);
sram_cell_6t_3 inst_cell_47_125 ( BL125, BLN125, WL47);
sram_cell_6t_3 inst_cell_47_124 ( BL124, BLN124, WL47);
sram_cell_6t_3 inst_cell_47_123 ( BL123, BLN123, WL47);
sram_cell_6t_3 inst_cell_47_122 ( BL122, BLN122, WL47);
sram_cell_6t_3 inst_cell_47_121 ( BL121, BLN121, WL47);
sram_cell_6t_3 inst_cell_47_120 ( BL120, BLN120, WL47);
sram_cell_6t_3 inst_cell_47_119 ( BL119, BLN119, WL47);
sram_cell_6t_3 inst_cell_47_118 ( BL118, BLN118, WL47);
sram_cell_6t_3 inst_cell_47_117 ( BL117, BLN117, WL47);
sram_cell_6t_3 inst_cell_47_116 ( BL116, BLN116, WL47);
sram_cell_6t_3 inst_cell_47_115 ( BL115, BLN115, WL47);
sram_cell_6t_3 inst_cell_47_114 ( BL114, BLN114, WL47);
sram_cell_6t_3 inst_cell_47_113 ( BL113, BLN113, WL47);
sram_cell_6t_3 inst_cell_47_112 ( BL112, BLN112, WL47);
sram_cell_6t_3 inst_cell_47_111 ( BL111, BLN111, WL47);
sram_cell_6t_3 inst_cell_47_110 ( BL110, BLN110, WL47);
sram_cell_6t_3 inst_cell_47_109 ( BL109, BLN109, WL47);
sram_cell_6t_3 inst_cell_47_108 ( BL108, BLN108, WL47);
sram_cell_6t_3 inst_cell_47_107 ( BL107, BLN107, WL47);
sram_cell_6t_3 inst_cell_47_106 ( BL106, BLN106, WL47);
sram_cell_6t_3 inst_cell_47_105 ( BL105, BLN105, WL47);
sram_cell_6t_3 inst_cell_47_104 ( BL104, BLN104, WL47);
sram_cell_6t_3 inst_cell_47_103 ( BL103, BLN103, WL47);
sram_cell_6t_3 inst_cell_47_102 ( BL102, BLN102, WL47);
sram_cell_6t_3 inst_cell_47_101 ( BL101, BLN101, WL47);
sram_cell_6t_3 inst_cell_47_100 ( BL100, BLN100, WL47);
sram_cell_6t_3 inst_cell_47_99 ( BL99, BLN99, WL47);
sram_cell_6t_3 inst_cell_47_98 ( BL98, BLN98, WL47);
sram_cell_6t_3 inst_cell_47_97 ( BL97, BLN97, WL47);
sram_cell_6t_3 inst_cell_47_96 ( BL96, BLN96, WL47);
sram_cell_6t_3 inst_cell_47_95 ( BL95, BLN95, WL47);
sram_cell_6t_3 inst_cell_47_94 ( BL94, BLN94, WL47);
sram_cell_6t_3 inst_cell_47_93 ( BL93, BLN93, WL47);
sram_cell_6t_3 inst_cell_47_92 ( BL92, BLN92, WL47);
sram_cell_6t_3 inst_cell_47_91 ( BL91, BLN91, WL47);
sram_cell_6t_3 inst_cell_47_90 ( BL90, BLN90, WL47);
sram_cell_6t_3 inst_cell_47_89 ( BL89, BLN89, WL47);
sram_cell_6t_3 inst_cell_47_88 ( BL88, BLN88, WL47);
sram_cell_6t_3 inst_cell_47_87 ( BL87, BLN87, WL47);
sram_cell_6t_3 inst_cell_47_86 ( BL86, BLN86, WL47);
sram_cell_6t_3 inst_cell_47_85 ( BL85, BLN85, WL47);
sram_cell_6t_3 inst_cell_47_84 ( BL84, BLN84, WL47);
sram_cell_6t_3 inst_cell_47_83 ( BL83, BLN83, WL47);
sram_cell_6t_3 inst_cell_47_82 ( BL82, BLN82, WL47);
sram_cell_6t_3 inst_cell_47_81 ( BL81, BLN81, WL47);
sram_cell_6t_3 inst_cell_47_80 ( BL80, BLN80, WL47);
sram_cell_6t_3 inst_cell_47_79 ( BL79, BLN79, WL47);
sram_cell_6t_3 inst_cell_47_78 ( BL78, BLN78, WL47);
sram_cell_6t_3 inst_cell_47_77 ( BL77, BLN77, WL47);
sram_cell_6t_3 inst_cell_47_76 ( BL76, BLN76, WL47);
sram_cell_6t_3 inst_cell_47_75 ( BL75, BLN75, WL47);
sram_cell_6t_3 inst_cell_47_74 ( BL74, BLN74, WL47);
sram_cell_6t_3 inst_cell_47_73 ( BL73, BLN73, WL47);
sram_cell_6t_3 inst_cell_47_72 ( BL72, BLN72, WL47);
sram_cell_6t_3 inst_cell_47_71 ( BL71, BLN71, WL47);
sram_cell_6t_3 inst_cell_47_70 ( BL70, BLN70, WL47);
sram_cell_6t_3 inst_cell_47_69 ( BL69, BLN69, WL47);
sram_cell_6t_3 inst_cell_47_68 ( BL68, BLN68, WL47);
sram_cell_6t_3 inst_cell_47_67 ( BL67, BLN67, WL47);
sram_cell_6t_3 inst_cell_47_66 ( BL66, BLN66, WL47);
sram_cell_6t_3 inst_cell_47_65 ( BL65, BLN65, WL47);
sram_cell_6t_3 inst_cell_47_64 ( BL64, BLN64, WL47);
sram_cell_6t_3 inst_cell_47_63 ( BL63, BLN63, WL47);
sram_cell_6t_3 inst_cell_47_62 ( BL62, BLN62, WL47);
sram_cell_6t_3 inst_cell_47_61 ( BL61, BLN61, WL47);
sram_cell_6t_3 inst_cell_47_60 ( BL60, BLN60, WL47);
sram_cell_6t_3 inst_cell_47_59 ( BL59, BLN59, WL47);
sram_cell_6t_3 inst_cell_47_58 ( BL58, BLN58, WL47);
sram_cell_6t_3 inst_cell_47_57 ( BL57, BLN57, WL47);
sram_cell_6t_3 inst_cell_47_56 ( BL56, BLN56, WL47);
sram_cell_6t_3 inst_cell_47_55 ( BL55, BLN55, WL47);
sram_cell_6t_3 inst_cell_47_54 ( BL54, BLN54, WL47);
sram_cell_6t_3 inst_cell_47_53 ( BL53, BLN53, WL47);
sram_cell_6t_3 inst_cell_47_52 ( BL52, BLN52, WL47);
sram_cell_6t_3 inst_cell_47_51 ( BL51, BLN51, WL47);
sram_cell_6t_3 inst_cell_47_50 ( BL50, BLN50, WL47);
sram_cell_6t_3 inst_cell_47_49 ( BL49, BLN49, WL47);
sram_cell_6t_3 inst_cell_47_48 ( BL48, BLN48, WL47);
sram_cell_6t_3 inst_cell_47_47 ( BL47, BLN47, WL47);
sram_cell_6t_3 inst_cell_47_46 ( BL46, BLN46, WL47);
sram_cell_6t_3 inst_cell_47_45 ( BL45, BLN45, WL47);
sram_cell_6t_3 inst_cell_47_44 ( BL44, BLN44, WL47);
sram_cell_6t_3 inst_cell_47_43 ( BL43, BLN43, WL47);
sram_cell_6t_3 inst_cell_47_42 ( BL42, BLN42, WL47);
sram_cell_6t_3 inst_cell_47_41 ( BL41, BLN41, WL47);
sram_cell_6t_3 inst_cell_47_40 ( BL40, BLN40, WL47);
sram_cell_6t_3 inst_cell_47_39 ( BL39, BLN39, WL47);
sram_cell_6t_3 inst_cell_47_38 ( BL38, BLN38, WL47);
sram_cell_6t_3 inst_cell_47_37 ( BL37, BLN37, WL47);
sram_cell_6t_3 inst_cell_47_36 ( BL36, BLN36, WL47);
sram_cell_6t_3 inst_cell_47_35 ( BL35, BLN35, WL47);
sram_cell_6t_3 inst_cell_47_34 ( BL34, BLN34, WL47);
sram_cell_6t_3 inst_cell_47_33 ( BL33, BLN33, WL47);
sram_cell_6t_3 inst_cell_47_32 ( BL32, BLN32, WL47);
sram_cell_6t_3 inst_cell_47_31 ( BL31, BLN31, WL47);
sram_cell_6t_3 inst_cell_47_30 ( BL30, BLN30, WL47);
sram_cell_6t_3 inst_cell_47_29 ( BL29, BLN29, WL47);
sram_cell_6t_3 inst_cell_47_28 ( BL28, BLN28, WL47);
sram_cell_6t_3 inst_cell_47_27 ( BL27, BLN27, WL47);
sram_cell_6t_3 inst_cell_47_26 ( BL26, BLN26, WL47);
sram_cell_6t_3 inst_cell_47_25 ( BL25, BLN25, WL47);
sram_cell_6t_3 inst_cell_47_24 ( BL24, BLN24, WL47);
sram_cell_6t_3 inst_cell_47_23 ( BL23, BLN23, WL47);
sram_cell_6t_3 inst_cell_47_22 ( BL22, BLN22, WL47);
sram_cell_6t_3 inst_cell_47_21 ( BL21, BLN21, WL47);
sram_cell_6t_3 inst_cell_47_20 ( BL20, BLN20, WL47);
sram_cell_6t_3 inst_cell_47_19 ( BL19, BLN19, WL47);
sram_cell_6t_3 inst_cell_47_18 ( BL18, BLN18, WL47);
sram_cell_6t_3 inst_cell_47_17 ( BL17, BLN17, WL47);
sram_cell_6t_3 inst_cell_47_16 ( BL16, BLN16, WL47);
sram_cell_6t_3 inst_cell_47_15 ( BL15, BLN15, WL47);
sram_cell_6t_3 inst_cell_47_14 ( BL14, BLN14, WL47);
sram_cell_6t_3 inst_cell_47_13 ( BL13, BLN13, WL47);
sram_cell_6t_3 inst_cell_47_12 ( BL12, BLN12, WL47);
sram_cell_6t_3 inst_cell_47_11 ( BL11, BLN11, WL47);
sram_cell_6t_3 inst_cell_47_10 ( BL10, BLN10, WL47);
sram_cell_6t_3 inst_cell_47_9 ( BL9, BLN9, WL47);
sram_cell_6t_3 inst_cell_47_8 ( BL8, BLN8, WL47);
sram_cell_6t_3 inst_cell_47_7 ( BL7, BLN7, WL47);
sram_cell_6t_3 inst_cell_47_6 ( BL6, BLN6, WL47);
sram_cell_6t_3 inst_cell_47_5 ( BL5, BLN5, WL47);
sram_cell_6t_3 inst_cell_47_4 ( BL4, BLN4, WL47);
sram_cell_6t_3 inst_cell_47_3 ( BL3, BLN3, WL47);
sram_cell_6t_3 inst_cell_47_2 ( BL2, BLN2, WL47);
sram_cell_6t_3 inst_cell_47_1 ( BL1, BLN1, WL47);
sram_cell_6t_3 inst_cell_47_0 ( BL0, BLN0, WL47);
sram_cell_6t_3 inst_cell_46_127 ( BL127, BLN127, WL46);
sram_cell_6t_3 inst_cell_46_126 ( BL126, BLN126, WL46);
sram_cell_6t_3 inst_cell_46_125 ( BL125, BLN125, WL46);
sram_cell_6t_3 inst_cell_46_124 ( BL124, BLN124, WL46);
sram_cell_6t_3 inst_cell_46_123 ( BL123, BLN123, WL46);
sram_cell_6t_3 inst_cell_46_122 ( BL122, BLN122, WL46);
sram_cell_6t_3 inst_cell_46_121 ( BL121, BLN121, WL46);
sram_cell_6t_3 inst_cell_46_120 ( BL120, BLN120, WL46);
sram_cell_6t_3 inst_cell_46_119 ( BL119, BLN119, WL46);
sram_cell_6t_3 inst_cell_46_118 ( BL118, BLN118, WL46);
sram_cell_6t_3 inst_cell_46_117 ( BL117, BLN117, WL46);
sram_cell_6t_3 inst_cell_46_116 ( BL116, BLN116, WL46);
sram_cell_6t_3 inst_cell_46_115 ( BL115, BLN115, WL46);
sram_cell_6t_3 inst_cell_46_114 ( BL114, BLN114, WL46);
sram_cell_6t_3 inst_cell_46_113 ( BL113, BLN113, WL46);
sram_cell_6t_3 inst_cell_46_112 ( BL112, BLN112, WL46);
sram_cell_6t_3 inst_cell_46_111 ( BL111, BLN111, WL46);
sram_cell_6t_3 inst_cell_46_110 ( BL110, BLN110, WL46);
sram_cell_6t_3 inst_cell_46_109 ( BL109, BLN109, WL46);
sram_cell_6t_3 inst_cell_46_108 ( BL108, BLN108, WL46);
sram_cell_6t_3 inst_cell_46_107 ( BL107, BLN107, WL46);
sram_cell_6t_3 inst_cell_46_106 ( BL106, BLN106, WL46);
sram_cell_6t_3 inst_cell_46_105 ( BL105, BLN105, WL46);
sram_cell_6t_3 inst_cell_46_104 ( BL104, BLN104, WL46);
sram_cell_6t_3 inst_cell_46_103 ( BL103, BLN103, WL46);
sram_cell_6t_3 inst_cell_46_102 ( BL102, BLN102, WL46);
sram_cell_6t_3 inst_cell_46_101 ( BL101, BLN101, WL46);
sram_cell_6t_3 inst_cell_46_100 ( BL100, BLN100, WL46);
sram_cell_6t_3 inst_cell_46_99 ( BL99, BLN99, WL46);
sram_cell_6t_3 inst_cell_46_98 ( BL98, BLN98, WL46);
sram_cell_6t_3 inst_cell_46_97 ( BL97, BLN97, WL46);
sram_cell_6t_3 inst_cell_46_96 ( BL96, BLN96, WL46);
sram_cell_6t_3 inst_cell_46_95 ( BL95, BLN95, WL46);
sram_cell_6t_3 inst_cell_46_94 ( BL94, BLN94, WL46);
sram_cell_6t_3 inst_cell_46_93 ( BL93, BLN93, WL46);
sram_cell_6t_3 inst_cell_46_92 ( BL92, BLN92, WL46);
sram_cell_6t_3 inst_cell_46_91 ( BL91, BLN91, WL46);
sram_cell_6t_3 inst_cell_46_90 ( BL90, BLN90, WL46);
sram_cell_6t_3 inst_cell_46_89 ( BL89, BLN89, WL46);
sram_cell_6t_3 inst_cell_46_88 ( BL88, BLN88, WL46);
sram_cell_6t_3 inst_cell_46_87 ( BL87, BLN87, WL46);
sram_cell_6t_3 inst_cell_46_86 ( BL86, BLN86, WL46);
sram_cell_6t_3 inst_cell_46_85 ( BL85, BLN85, WL46);
sram_cell_6t_3 inst_cell_46_84 ( BL84, BLN84, WL46);
sram_cell_6t_3 inst_cell_46_83 ( BL83, BLN83, WL46);
sram_cell_6t_3 inst_cell_46_82 ( BL82, BLN82, WL46);
sram_cell_6t_3 inst_cell_46_81 ( BL81, BLN81, WL46);
sram_cell_6t_3 inst_cell_46_80 ( BL80, BLN80, WL46);
sram_cell_6t_3 inst_cell_46_79 ( BL79, BLN79, WL46);
sram_cell_6t_3 inst_cell_46_78 ( BL78, BLN78, WL46);
sram_cell_6t_3 inst_cell_46_77 ( BL77, BLN77, WL46);
sram_cell_6t_3 inst_cell_46_76 ( BL76, BLN76, WL46);
sram_cell_6t_3 inst_cell_46_75 ( BL75, BLN75, WL46);
sram_cell_6t_3 inst_cell_46_74 ( BL74, BLN74, WL46);
sram_cell_6t_3 inst_cell_46_73 ( BL73, BLN73, WL46);
sram_cell_6t_3 inst_cell_46_72 ( BL72, BLN72, WL46);
sram_cell_6t_3 inst_cell_46_71 ( BL71, BLN71, WL46);
sram_cell_6t_3 inst_cell_46_70 ( BL70, BLN70, WL46);
sram_cell_6t_3 inst_cell_46_69 ( BL69, BLN69, WL46);
sram_cell_6t_3 inst_cell_46_68 ( BL68, BLN68, WL46);
sram_cell_6t_3 inst_cell_46_67 ( BL67, BLN67, WL46);
sram_cell_6t_3 inst_cell_46_66 ( BL66, BLN66, WL46);
sram_cell_6t_3 inst_cell_46_65 ( BL65, BLN65, WL46);
sram_cell_6t_3 inst_cell_46_64 ( BL64, BLN64, WL46);
sram_cell_6t_3 inst_cell_46_63 ( BL63, BLN63, WL46);
sram_cell_6t_3 inst_cell_46_62 ( BL62, BLN62, WL46);
sram_cell_6t_3 inst_cell_46_61 ( BL61, BLN61, WL46);
sram_cell_6t_3 inst_cell_46_60 ( BL60, BLN60, WL46);
sram_cell_6t_3 inst_cell_46_59 ( BL59, BLN59, WL46);
sram_cell_6t_3 inst_cell_46_58 ( BL58, BLN58, WL46);
sram_cell_6t_3 inst_cell_46_57 ( BL57, BLN57, WL46);
sram_cell_6t_3 inst_cell_46_56 ( BL56, BLN56, WL46);
sram_cell_6t_3 inst_cell_46_55 ( BL55, BLN55, WL46);
sram_cell_6t_3 inst_cell_46_54 ( BL54, BLN54, WL46);
sram_cell_6t_3 inst_cell_46_53 ( BL53, BLN53, WL46);
sram_cell_6t_3 inst_cell_46_52 ( BL52, BLN52, WL46);
sram_cell_6t_3 inst_cell_46_51 ( BL51, BLN51, WL46);
sram_cell_6t_3 inst_cell_46_50 ( BL50, BLN50, WL46);
sram_cell_6t_3 inst_cell_46_49 ( BL49, BLN49, WL46);
sram_cell_6t_3 inst_cell_46_48 ( BL48, BLN48, WL46);
sram_cell_6t_3 inst_cell_46_47 ( BL47, BLN47, WL46);
sram_cell_6t_3 inst_cell_46_46 ( BL46, BLN46, WL46);
sram_cell_6t_3 inst_cell_46_45 ( BL45, BLN45, WL46);
sram_cell_6t_3 inst_cell_46_44 ( BL44, BLN44, WL46);
sram_cell_6t_3 inst_cell_46_43 ( BL43, BLN43, WL46);
sram_cell_6t_3 inst_cell_46_42 ( BL42, BLN42, WL46);
sram_cell_6t_3 inst_cell_46_41 ( BL41, BLN41, WL46);
sram_cell_6t_3 inst_cell_46_40 ( BL40, BLN40, WL46);
sram_cell_6t_3 inst_cell_46_39 ( BL39, BLN39, WL46);
sram_cell_6t_3 inst_cell_46_38 ( BL38, BLN38, WL46);
sram_cell_6t_3 inst_cell_46_37 ( BL37, BLN37, WL46);
sram_cell_6t_3 inst_cell_46_36 ( BL36, BLN36, WL46);
sram_cell_6t_3 inst_cell_46_35 ( BL35, BLN35, WL46);
sram_cell_6t_3 inst_cell_46_34 ( BL34, BLN34, WL46);
sram_cell_6t_3 inst_cell_46_33 ( BL33, BLN33, WL46);
sram_cell_6t_3 inst_cell_46_32 ( BL32, BLN32, WL46);
sram_cell_6t_3 inst_cell_46_31 ( BL31, BLN31, WL46);
sram_cell_6t_3 inst_cell_46_30 ( BL30, BLN30, WL46);
sram_cell_6t_3 inst_cell_46_29 ( BL29, BLN29, WL46);
sram_cell_6t_3 inst_cell_46_28 ( BL28, BLN28, WL46);
sram_cell_6t_3 inst_cell_46_27 ( BL27, BLN27, WL46);
sram_cell_6t_3 inst_cell_46_26 ( BL26, BLN26, WL46);
sram_cell_6t_3 inst_cell_46_25 ( BL25, BLN25, WL46);
sram_cell_6t_3 inst_cell_46_24 ( BL24, BLN24, WL46);
sram_cell_6t_3 inst_cell_46_23 ( BL23, BLN23, WL46);
sram_cell_6t_3 inst_cell_46_22 ( BL22, BLN22, WL46);
sram_cell_6t_3 inst_cell_46_21 ( BL21, BLN21, WL46);
sram_cell_6t_3 inst_cell_46_20 ( BL20, BLN20, WL46);
sram_cell_6t_3 inst_cell_46_19 ( BL19, BLN19, WL46);
sram_cell_6t_3 inst_cell_46_18 ( BL18, BLN18, WL46);
sram_cell_6t_3 inst_cell_46_17 ( BL17, BLN17, WL46);
sram_cell_6t_3 inst_cell_46_16 ( BL16, BLN16, WL46);
sram_cell_6t_3 inst_cell_46_15 ( BL15, BLN15, WL46);
sram_cell_6t_3 inst_cell_46_14 ( BL14, BLN14, WL46);
sram_cell_6t_3 inst_cell_46_13 ( BL13, BLN13, WL46);
sram_cell_6t_3 inst_cell_46_12 ( BL12, BLN12, WL46);
sram_cell_6t_3 inst_cell_46_11 ( BL11, BLN11, WL46);
sram_cell_6t_3 inst_cell_46_10 ( BL10, BLN10, WL46);
sram_cell_6t_3 inst_cell_46_9 ( BL9, BLN9, WL46);
sram_cell_6t_3 inst_cell_46_8 ( BL8, BLN8, WL46);
sram_cell_6t_3 inst_cell_46_7 ( BL7, BLN7, WL46);
sram_cell_6t_3 inst_cell_46_6 ( BL6, BLN6, WL46);
sram_cell_6t_3 inst_cell_46_5 ( BL5, BLN5, WL46);
sram_cell_6t_3 inst_cell_46_4 ( BL4, BLN4, WL46);
sram_cell_6t_3 inst_cell_46_3 ( BL3, BLN3, WL46);
sram_cell_6t_3 inst_cell_46_2 ( BL2, BLN2, WL46);
sram_cell_6t_3 inst_cell_46_1 ( BL1, BLN1, WL46);
sram_cell_6t_3 inst_cell_46_0 ( BL0, BLN0, WL46);
sram_cell_6t_3 inst_cell_45_127 ( BL127, BLN127, WL45);
sram_cell_6t_3 inst_cell_45_126 ( BL126, BLN126, WL45);
sram_cell_6t_3 inst_cell_45_125 ( BL125, BLN125, WL45);
sram_cell_6t_3 inst_cell_45_124 ( BL124, BLN124, WL45);
sram_cell_6t_3 inst_cell_45_123 ( BL123, BLN123, WL45);
sram_cell_6t_3 inst_cell_45_122 ( BL122, BLN122, WL45);
sram_cell_6t_3 inst_cell_45_121 ( BL121, BLN121, WL45);
sram_cell_6t_3 inst_cell_45_120 ( BL120, BLN120, WL45);
sram_cell_6t_3 inst_cell_45_119 ( BL119, BLN119, WL45);
sram_cell_6t_3 inst_cell_45_118 ( BL118, BLN118, WL45);
sram_cell_6t_3 inst_cell_45_117 ( BL117, BLN117, WL45);
sram_cell_6t_3 inst_cell_45_116 ( BL116, BLN116, WL45);
sram_cell_6t_3 inst_cell_45_115 ( BL115, BLN115, WL45);
sram_cell_6t_3 inst_cell_45_114 ( BL114, BLN114, WL45);
sram_cell_6t_3 inst_cell_45_113 ( BL113, BLN113, WL45);
sram_cell_6t_3 inst_cell_45_112 ( BL112, BLN112, WL45);
sram_cell_6t_3 inst_cell_45_111 ( BL111, BLN111, WL45);
sram_cell_6t_3 inst_cell_45_110 ( BL110, BLN110, WL45);
sram_cell_6t_3 inst_cell_45_109 ( BL109, BLN109, WL45);
sram_cell_6t_3 inst_cell_45_108 ( BL108, BLN108, WL45);
sram_cell_6t_3 inst_cell_45_107 ( BL107, BLN107, WL45);
sram_cell_6t_3 inst_cell_45_106 ( BL106, BLN106, WL45);
sram_cell_6t_3 inst_cell_45_105 ( BL105, BLN105, WL45);
sram_cell_6t_3 inst_cell_45_104 ( BL104, BLN104, WL45);
sram_cell_6t_3 inst_cell_45_103 ( BL103, BLN103, WL45);
sram_cell_6t_3 inst_cell_45_102 ( BL102, BLN102, WL45);
sram_cell_6t_3 inst_cell_45_101 ( BL101, BLN101, WL45);
sram_cell_6t_3 inst_cell_45_100 ( BL100, BLN100, WL45);
sram_cell_6t_3 inst_cell_45_99 ( BL99, BLN99, WL45);
sram_cell_6t_3 inst_cell_45_98 ( BL98, BLN98, WL45);
sram_cell_6t_3 inst_cell_45_97 ( BL97, BLN97, WL45);
sram_cell_6t_3 inst_cell_45_96 ( BL96, BLN96, WL45);
sram_cell_6t_3 inst_cell_45_95 ( BL95, BLN95, WL45);
sram_cell_6t_3 inst_cell_45_94 ( BL94, BLN94, WL45);
sram_cell_6t_3 inst_cell_45_93 ( BL93, BLN93, WL45);
sram_cell_6t_3 inst_cell_45_92 ( BL92, BLN92, WL45);
sram_cell_6t_3 inst_cell_45_91 ( BL91, BLN91, WL45);
sram_cell_6t_3 inst_cell_45_90 ( BL90, BLN90, WL45);
sram_cell_6t_3 inst_cell_45_89 ( BL89, BLN89, WL45);
sram_cell_6t_3 inst_cell_45_88 ( BL88, BLN88, WL45);
sram_cell_6t_3 inst_cell_45_87 ( BL87, BLN87, WL45);
sram_cell_6t_3 inst_cell_45_86 ( BL86, BLN86, WL45);
sram_cell_6t_3 inst_cell_45_85 ( BL85, BLN85, WL45);
sram_cell_6t_3 inst_cell_45_84 ( BL84, BLN84, WL45);
sram_cell_6t_3 inst_cell_45_83 ( BL83, BLN83, WL45);
sram_cell_6t_3 inst_cell_45_82 ( BL82, BLN82, WL45);
sram_cell_6t_3 inst_cell_45_81 ( BL81, BLN81, WL45);
sram_cell_6t_3 inst_cell_45_80 ( BL80, BLN80, WL45);
sram_cell_6t_3 inst_cell_45_79 ( BL79, BLN79, WL45);
sram_cell_6t_3 inst_cell_45_78 ( BL78, BLN78, WL45);
sram_cell_6t_3 inst_cell_45_77 ( BL77, BLN77, WL45);
sram_cell_6t_3 inst_cell_45_76 ( BL76, BLN76, WL45);
sram_cell_6t_3 inst_cell_45_75 ( BL75, BLN75, WL45);
sram_cell_6t_3 inst_cell_45_74 ( BL74, BLN74, WL45);
sram_cell_6t_3 inst_cell_45_73 ( BL73, BLN73, WL45);
sram_cell_6t_3 inst_cell_45_72 ( BL72, BLN72, WL45);
sram_cell_6t_3 inst_cell_45_71 ( BL71, BLN71, WL45);
sram_cell_6t_3 inst_cell_45_70 ( BL70, BLN70, WL45);
sram_cell_6t_3 inst_cell_45_69 ( BL69, BLN69, WL45);
sram_cell_6t_3 inst_cell_45_68 ( BL68, BLN68, WL45);
sram_cell_6t_3 inst_cell_45_67 ( BL67, BLN67, WL45);
sram_cell_6t_3 inst_cell_45_66 ( BL66, BLN66, WL45);
sram_cell_6t_3 inst_cell_45_65 ( BL65, BLN65, WL45);
sram_cell_6t_3 inst_cell_45_64 ( BL64, BLN64, WL45);
sram_cell_6t_3 inst_cell_45_63 ( BL63, BLN63, WL45);
sram_cell_6t_3 inst_cell_45_62 ( BL62, BLN62, WL45);
sram_cell_6t_3 inst_cell_45_61 ( BL61, BLN61, WL45);
sram_cell_6t_3 inst_cell_45_60 ( BL60, BLN60, WL45);
sram_cell_6t_3 inst_cell_45_59 ( BL59, BLN59, WL45);
sram_cell_6t_3 inst_cell_45_58 ( BL58, BLN58, WL45);
sram_cell_6t_3 inst_cell_45_57 ( BL57, BLN57, WL45);
sram_cell_6t_3 inst_cell_45_56 ( BL56, BLN56, WL45);
sram_cell_6t_3 inst_cell_45_55 ( BL55, BLN55, WL45);
sram_cell_6t_3 inst_cell_45_54 ( BL54, BLN54, WL45);
sram_cell_6t_3 inst_cell_45_53 ( BL53, BLN53, WL45);
sram_cell_6t_3 inst_cell_45_52 ( BL52, BLN52, WL45);
sram_cell_6t_3 inst_cell_45_51 ( BL51, BLN51, WL45);
sram_cell_6t_3 inst_cell_45_50 ( BL50, BLN50, WL45);
sram_cell_6t_3 inst_cell_45_49 ( BL49, BLN49, WL45);
sram_cell_6t_3 inst_cell_45_48 ( BL48, BLN48, WL45);
sram_cell_6t_3 inst_cell_45_47 ( BL47, BLN47, WL45);
sram_cell_6t_3 inst_cell_45_46 ( BL46, BLN46, WL45);
sram_cell_6t_3 inst_cell_45_45 ( BL45, BLN45, WL45);
sram_cell_6t_3 inst_cell_45_44 ( BL44, BLN44, WL45);
sram_cell_6t_3 inst_cell_45_43 ( BL43, BLN43, WL45);
sram_cell_6t_3 inst_cell_45_42 ( BL42, BLN42, WL45);
sram_cell_6t_3 inst_cell_45_41 ( BL41, BLN41, WL45);
sram_cell_6t_3 inst_cell_45_40 ( BL40, BLN40, WL45);
sram_cell_6t_3 inst_cell_45_39 ( BL39, BLN39, WL45);
sram_cell_6t_3 inst_cell_45_38 ( BL38, BLN38, WL45);
sram_cell_6t_3 inst_cell_45_37 ( BL37, BLN37, WL45);
sram_cell_6t_3 inst_cell_45_36 ( BL36, BLN36, WL45);
sram_cell_6t_3 inst_cell_45_35 ( BL35, BLN35, WL45);
sram_cell_6t_3 inst_cell_45_34 ( BL34, BLN34, WL45);
sram_cell_6t_3 inst_cell_45_33 ( BL33, BLN33, WL45);
sram_cell_6t_3 inst_cell_45_32 ( BL32, BLN32, WL45);
sram_cell_6t_3 inst_cell_45_31 ( BL31, BLN31, WL45);
sram_cell_6t_3 inst_cell_45_30 ( BL30, BLN30, WL45);
sram_cell_6t_3 inst_cell_45_29 ( BL29, BLN29, WL45);
sram_cell_6t_3 inst_cell_45_28 ( BL28, BLN28, WL45);
sram_cell_6t_3 inst_cell_45_27 ( BL27, BLN27, WL45);
sram_cell_6t_3 inst_cell_45_26 ( BL26, BLN26, WL45);
sram_cell_6t_3 inst_cell_45_25 ( BL25, BLN25, WL45);
sram_cell_6t_3 inst_cell_45_24 ( BL24, BLN24, WL45);
sram_cell_6t_3 inst_cell_45_23 ( BL23, BLN23, WL45);
sram_cell_6t_3 inst_cell_45_22 ( BL22, BLN22, WL45);
sram_cell_6t_3 inst_cell_45_21 ( BL21, BLN21, WL45);
sram_cell_6t_3 inst_cell_45_20 ( BL20, BLN20, WL45);
sram_cell_6t_3 inst_cell_45_19 ( BL19, BLN19, WL45);
sram_cell_6t_3 inst_cell_45_18 ( BL18, BLN18, WL45);
sram_cell_6t_3 inst_cell_45_17 ( BL17, BLN17, WL45);
sram_cell_6t_3 inst_cell_45_16 ( BL16, BLN16, WL45);
sram_cell_6t_3 inst_cell_45_15 ( BL15, BLN15, WL45);
sram_cell_6t_3 inst_cell_45_14 ( BL14, BLN14, WL45);
sram_cell_6t_3 inst_cell_45_13 ( BL13, BLN13, WL45);
sram_cell_6t_3 inst_cell_45_12 ( BL12, BLN12, WL45);
sram_cell_6t_3 inst_cell_45_11 ( BL11, BLN11, WL45);
sram_cell_6t_3 inst_cell_45_10 ( BL10, BLN10, WL45);
sram_cell_6t_3 inst_cell_45_9 ( BL9, BLN9, WL45);
sram_cell_6t_3 inst_cell_45_8 ( BL8, BLN8, WL45);
sram_cell_6t_3 inst_cell_45_7 ( BL7, BLN7, WL45);
sram_cell_6t_3 inst_cell_45_6 ( BL6, BLN6, WL45);
sram_cell_6t_3 inst_cell_45_5 ( BL5, BLN5, WL45);
sram_cell_6t_3 inst_cell_45_4 ( BL4, BLN4, WL45);
sram_cell_6t_3 inst_cell_45_3 ( BL3, BLN3, WL45);
sram_cell_6t_3 inst_cell_45_2 ( BL2, BLN2, WL45);
sram_cell_6t_3 inst_cell_45_1 ( BL1, BLN1, WL45);
sram_cell_6t_3 inst_cell_45_0 ( BL0, BLN0, WL45);
sram_cell_6t_3 inst_cell_44_127 ( BL127, BLN127, WL44);
sram_cell_6t_3 inst_cell_44_126 ( BL126, BLN126, WL44);
sram_cell_6t_3 inst_cell_44_125 ( BL125, BLN125, WL44);
sram_cell_6t_3 inst_cell_44_124 ( BL124, BLN124, WL44);
sram_cell_6t_3 inst_cell_44_123 ( BL123, BLN123, WL44);
sram_cell_6t_3 inst_cell_44_122 ( BL122, BLN122, WL44);
sram_cell_6t_3 inst_cell_44_121 ( BL121, BLN121, WL44);
sram_cell_6t_3 inst_cell_44_120 ( BL120, BLN120, WL44);
sram_cell_6t_3 inst_cell_44_119 ( BL119, BLN119, WL44);
sram_cell_6t_3 inst_cell_44_118 ( BL118, BLN118, WL44);
sram_cell_6t_3 inst_cell_44_117 ( BL117, BLN117, WL44);
sram_cell_6t_3 inst_cell_44_116 ( BL116, BLN116, WL44);
sram_cell_6t_3 inst_cell_44_115 ( BL115, BLN115, WL44);
sram_cell_6t_3 inst_cell_44_114 ( BL114, BLN114, WL44);
sram_cell_6t_3 inst_cell_44_113 ( BL113, BLN113, WL44);
sram_cell_6t_3 inst_cell_44_112 ( BL112, BLN112, WL44);
sram_cell_6t_3 inst_cell_44_111 ( BL111, BLN111, WL44);
sram_cell_6t_3 inst_cell_44_110 ( BL110, BLN110, WL44);
sram_cell_6t_3 inst_cell_44_109 ( BL109, BLN109, WL44);
sram_cell_6t_3 inst_cell_44_108 ( BL108, BLN108, WL44);
sram_cell_6t_3 inst_cell_44_107 ( BL107, BLN107, WL44);
sram_cell_6t_3 inst_cell_44_106 ( BL106, BLN106, WL44);
sram_cell_6t_3 inst_cell_44_105 ( BL105, BLN105, WL44);
sram_cell_6t_3 inst_cell_44_104 ( BL104, BLN104, WL44);
sram_cell_6t_3 inst_cell_44_103 ( BL103, BLN103, WL44);
sram_cell_6t_3 inst_cell_44_102 ( BL102, BLN102, WL44);
sram_cell_6t_3 inst_cell_44_101 ( BL101, BLN101, WL44);
sram_cell_6t_3 inst_cell_44_100 ( BL100, BLN100, WL44);
sram_cell_6t_3 inst_cell_44_99 ( BL99, BLN99, WL44);
sram_cell_6t_3 inst_cell_44_98 ( BL98, BLN98, WL44);
sram_cell_6t_3 inst_cell_44_97 ( BL97, BLN97, WL44);
sram_cell_6t_3 inst_cell_44_96 ( BL96, BLN96, WL44);
sram_cell_6t_3 inst_cell_44_95 ( BL95, BLN95, WL44);
sram_cell_6t_3 inst_cell_44_94 ( BL94, BLN94, WL44);
sram_cell_6t_3 inst_cell_44_93 ( BL93, BLN93, WL44);
sram_cell_6t_3 inst_cell_44_92 ( BL92, BLN92, WL44);
sram_cell_6t_3 inst_cell_44_91 ( BL91, BLN91, WL44);
sram_cell_6t_3 inst_cell_44_90 ( BL90, BLN90, WL44);
sram_cell_6t_3 inst_cell_44_89 ( BL89, BLN89, WL44);
sram_cell_6t_3 inst_cell_44_88 ( BL88, BLN88, WL44);
sram_cell_6t_3 inst_cell_44_87 ( BL87, BLN87, WL44);
sram_cell_6t_3 inst_cell_44_86 ( BL86, BLN86, WL44);
sram_cell_6t_3 inst_cell_44_85 ( BL85, BLN85, WL44);
sram_cell_6t_3 inst_cell_44_84 ( BL84, BLN84, WL44);
sram_cell_6t_3 inst_cell_44_83 ( BL83, BLN83, WL44);
sram_cell_6t_3 inst_cell_44_82 ( BL82, BLN82, WL44);
sram_cell_6t_3 inst_cell_44_81 ( BL81, BLN81, WL44);
sram_cell_6t_3 inst_cell_44_80 ( BL80, BLN80, WL44);
sram_cell_6t_3 inst_cell_44_79 ( BL79, BLN79, WL44);
sram_cell_6t_3 inst_cell_44_78 ( BL78, BLN78, WL44);
sram_cell_6t_3 inst_cell_44_77 ( BL77, BLN77, WL44);
sram_cell_6t_3 inst_cell_44_76 ( BL76, BLN76, WL44);
sram_cell_6t_3 inst_cell_44_75 ( BL75, BLN75, WL44);
sram_cell_6t_3 inst_cell_44_74 ( BL74, BLN74, WL44);
sram_cell_6t_3 inst_cell_44_73 ( BL73, BLN73, WL44);
sram_cell_6t_3 inst_cell_44_72 ( BL72, BLN72, WL44);
sram_cell_6t_3 inst_cell_44_71 ( BL71, BLN71, WL44);
sram_cell_6t_3 inst_cell_44_70 ( BL70, BLN70, WL44);
sram_cell_6t_3 inst_cell_44_69 ( BL69, BLN69, WL44);
sram_cell_6t_3 inst_cell_44_68 ( BL68, BLN68, WL44);
sram_cell_6t_3 inst_cell_44_67 ( BL67, BLN67, WL44);
sram_cell_6t_3 inst_cell_44_66 ( BL66, BLN66, WL44);
sram_cell_6t_3 inst_cell_44_65 ( BL65, BLN65, WL44);
sram_cell_6t_3 inst_cell_44_64 ( BL64, BLN64, WL44);
sram_cell_6t_3 inst_cell_44_63 ( BL63, BLN63, WL44);
sram_cell_6t_3 inst_cell_44_62 ( BL62, BLN62, WL44);
sram_cell_6t_3 inst_cell_44_61 ( BL61, BLN61, WL44);
sram_cell_6t_3 inst_cell_44_60 ( BL60, BLN60, WL44);
sram_cell_6t_3 inst_cell_44_59 ( BL59, BLN59, WL44);
sram_cell_6t_3 inst_cell_44_58 ( BL58, BLN58, WL44);
sram_cell_6t_3 inst_cell_44_57 ( BL57, BLN57, WL44);
sram_cell_6t_3 inst_cell_44_56 ( BL56, BLN56, WL44);
sram_cell_6t_3 inst_cell_44_55 ( BL55, BLN55, WL44);
sram_cell_6t_3 inst_cell_44_54 ( BL54, BLN54, WL44);
sram_cell_6t_3 inst_cell_44_53 ( BL53, BLN53, WL44);
sram_cell_6t_3 inst_cell_44_52 ( BL52, BLN52, WL44);
sram_cell_6t_3 inst_cell_44_51 ( BL51, BLN51, WL44);
sram_cell_6t_3 inst_cell_44_50 ( BL50, BLN50, WL44);
sram_cell_6t_3 inst_cell_44_49 ( BL49, BLN49, WL44);
sram_cell_6t_3 inst_cell_44_48 ( BL48, BLN48, WL44);
sram_cell_6t_3 inst_cell_44_47 ( BL47, BLN47, WL44);
sram_cell_6t_3 inst_cell_44_46 ( BL46, BLN46, WL44);
sram_cell_6t_3 inst_cell_44_45 ( BL45, BLN45, WL44);
sram_cell_6t_3 inst_cell_44_44 ( BL44, BLN44, WL44);
sram_cell_6t_3 inst_cell_44_43 ( BL43, BLN43, WL44);
sram_cell_6t_3 inst_cell_44_42 ( BL42, BLN42, WL44);
sram_cell_6t_3 inst_cell_44_41 ( BL41, BLN41, WL44);
sram_cell_6t_3 inst_cell_44_40 ( BL40, BLN40, WL44);
sram_cell_6t_3 inst_cell_44_39 ( BL39, BLN39, WL44);
sram_cell_6t_3 inst_cell_44_38 ( BL38, BLN38, WL44);
sram_cell_6t_3 inst_cell_44_37 ( BL37, BLN37, WL44);
sram_cell_6t_3 inst_cell_44_36 ( BL36, BLN36, WL44);
sram_cell_6t_3 inst_cell_44_35 ( BL35, BLN35, WL44);
sram_cell_6t_3 inst_cell_44_34 ( BL34, BLN34, WL44);
sram_cell_6t_3 inst_cell_44_33 ( BL33, BLN33, WL44);
sram_cell_6t_3 inst_cell_44_32 ( BL32, BLN32, WL44);
sram_cell_6t_3 inst_cell_44_31 ( BL31, BLN31, WL44);
sram_cell_6t_3 inst_cell_44_30 ( BL30, BLN30, WL44);
sram_cell_6t_3 inst_cell_44_29 ( BL29, BLN29, WL44);
sram_cell_6t_3 inst_cell_44_28 ( BL28, BLN28, WL44);
sram_cell_6t_3 inst_cell_44_27 ( BL27, BLN27, WL44);
sram_cell_6t_3 inst_cell_44_26 ( BL26, BLN26, WL44);
sram_cell_6t_3 inst_cell_44_25 ( BL25, BLN25, WL44);
sram_cell_6t_3 inst_cell_44_24 ( BL24, BLN24, WL44);
sram_cell_6t_3 inst_cell_44_23 ( BL23, BLN23, WL44);
sram_cell_6t_3 inst_cell_44_22 ( BL22, BLN22, WL44);
sram_cell_6t_3 inst_cell_44_21 ( BL21, BLN21, WL44);
sram_cell_6t_3 inst_cell_44_20 ( BL20, BLN20, WL44);
sram_cell_6t_3 inst_cell_44_19 ( BL19, BLN19, WL44);
sram_cell_6t_3 inst_cell_44_18 ( BL18, BLN18, WL44);
sram_cell_6t_3 inst_cell_44_17 ( BL17, BLN17, WL44);
sram_cell_6t_3 inst_cell_44_16 ( BL16, BLN16, WL44);
sram_cell_6t_3 inst_cell_44_15 ( BL15, BLN15, WL44);
sram_cell_6t_3 inst_cell_44_14 ( BL14, BLN14, WL44);
sram_cell_6t_3 inst_cell_44_13 ( BL13, BLN13, WL44);
sram_cell_6t_3 inst_cell_44_12 ( BL12, BLN12, WL44);
sram_cell_6t_3 inst_cell_44_11 ( BL11, BLN11, WL44);
sram_cell_6t_3 inst_cell_44_10 ( BL10, BLN10, WL44);
sram_cell_6t_3 inst_cell_44_9 ( BL9, BLN9, WL44);
sram_cell_6t_3 inst_cell_44_8 ( BL8, BLN8, WL44);
sram_cell_6t_3 inst_cell_44_7 ( BL7, BLN7, WL44);
sram_cell_6t_3 inst_cell_44_6 ( BL6, BLN6, WL44);
sram_cell_6t_3 inst_cell_44_5 ( BL5, BLN5, WL44);
sram_cell_6t_3 inst_cell_44_4 ( BL4, BLN4, WL44);
sram_cell_6t_3 inst_cell_44_3 ( BL3, BLN3, WL44);
sram_cell_6t_3 inst_cell_44_2 ( BL2, BLN2, WL44);
sram_cell_6t_3 inst_cell_44_1 ( BL1, BLN1, WL44);
sram_cell_6t_3 inst_cell_44_0 ( BL0, BLN0, WL44);
sram_cell_6t_3 inst_cell_43_127 ( BL127, BLN127, WL43);
sram_cell_6t_3 inst_cell_43_126 ( BL126, BLN126, WL43);
sram_cell_6t_3 inst_cell_43_125 ( BL125, BLN125, WL43);
sram_cell_6t_3 inst_cell_43_124 ( BL124, BLN124, WL43);
sram_cell_6t_3 inst_cell_43_123 ( BL123, BLN123, WL43);
sram_cell_6t_3 inst_cell_43_122 ( BL122, BLN122, WL43);
sram_cell_6t_3 inst_cell_43_121 ( BL121, BLN121, WL43);
sram_cell_6t_3 inst_cell_43_120 ( BL120, BLN120, WL43);
sram_cell_6t_3 inst_cell_43_119 ( BL119, BLN119, WL43);
sram_cell_6t_3 inst_cell_43_118 ( BL118, BLN118, WL43);
sram_cell_6t_3 inst_cell_43_117 ( BL117, BLN117, WL43);
sram_cell_6t_3 inst_cell_43_116 ( BL116, BLN116, WL43);
sram_cell_6t_3 inst_cell_43_115 ( BL115, BLN115, WL43);
sram_cell_6t_3 inst_cell_43_114 ( BL114, BLN114, WL43);
sram_cell_6t_3 inst_cell_43_113 ( BL113, BLN113, WL43);
sram_cell_6t_3 inst_cell_43_112 ( BL112, BLN112, WL43);
sram_cell_6t_3 inst_cell_43_111 ( BL111, BLN111, WL43);
sram_cell_6t_3 inst_cell_43_110 ( BL110, BLN110, WL43);
sram_cell_6t_3 inst_cell_43_109 ( BL109, BLN109, WL43);
sram_cell_6t_3 inst_cell_43_108 ( BL108, BLN108, WL43);
sram_cell_6t_3 inst_cell_43_107 ( BL107, BLN107, WL43);
sram_cell_6t_3 inst_cell_43_106 ( BL106, BLN106, WL43);
sram_cell_6t_3 inst_cell_43_105 ( BL105, BLN105, WL43);
sram_cell_6t_3 inst_cell_43_104 ( BL104, BLN104, WL43);
sram_cell_6t_3 inst_cell_43_103 ( BL103, BLN103, WL43);
sram_cell_6t_3 inst_cell_43_102 ( BL102, BLN102, WL43);
sram_cell_6t_3 inst_cell_43_101 ( BL101, BLN101, WL43);
sram_cell_6t_3 inst_cell_43_100 ( BL100, BLN100, WL43);
sram_cell_6t_3 inst_cell_43_99 ( BL99, BLN99, WL43);
sram_cell_6t_3 inst_cell_43_98 ( BL98, BLN98, WL43);
sram_cell_6t_3 inst_cell_43_97 ( BL97, BLN97, WL43);
sram_cell_6t_3 inst_cell_43_96 ( BL96, BLN96, WL43);
sram_cell_6t_3 inst_cell_43_95 ( BL95, BLN95, WL43);
sram_cell_6t_3 inst_cell_43_94 ( BL94, BLN94, WL43);
sram_cell_6t_3 inst_cell_43_93 ( BL93, BLN93, WL43);
sram_cell_6t_3 inst_cell_43_92 ( BL92, BLN92, WL43);
sram_cell_6t_3 inst_cell_43_91 ( BL91, BLN91, WL43);
sram_cell_6t_3 inst_cell_43_90 ( BL90, BLN90, WL43);
sram_cell_6t_3 inst_cell_43_89 ( BL89, BLN89, WL43);
sram_cell_6t_3 inst_cell_43_88 ( BL88, BLN88, WL43);
sram_cell_6t_3 inst_cell_43_87 ( BL87, BLN87, WL43);
sram_cell_6t_3 inst_cell_43_86 ( BL86, BLN86, WL43);
sram_cell_6t_3 inst_cell_43_85 ( BL85, BLN85, WL43);
sram_cell_6t_3 inst_cell_43_84 ( BL84, BLN84, WL43);
sram_cell_6t_3 inst_cell_43_83 ( BL83, BLN83, WL43);
sram_cell_6t_3 inst_cell_43_82 ( BL82, BLN82, WL43);
sram_cell_6t_3 inst_cell_43_81 ( BL81, BLN81, WL43);
sram_cell_6t_3 inst_cell_43_80 ( BL80, BLN80, WL43);
sram_cell_6t_3 inst_cell_43_79 ( BL79, BLN79, WL43);
sram_cell_6t_3 inst_cell_43_78 ( BL78, BLN78, WL43);
sram_cell_6t_3 inst_cell_43_77 ( BL77, BLN77, WL43);
sram_cell_6t_3 inst_cell_43_76 ( BL76, BLN76, WL43);
sram_cell_6t_3 inst_cell_43_75 ( BL75, BLN75, WL43);
sram_cell_6t_3 inst_cell_43_74 ( BL74, BLN74, WL43);
sram_cell_6t_3 inst_cell_43_73 ( BL73, BLN73, WL43);
sram_cell_6t_3 inst_cell_43_72 ( BL72, BLN72, WL43);
sram_cell_6t_3 inst_cell_43_71 ( BL71, BLN71, WL43);
sram_cell_6t_3 inst_cell_43_70 ( BL70, BLN70, WL43);
sram_cell_6t_3 inst_cell_43_69 ( BL69, BLN69, WL43);
sram_cell_6t_3 inst_cell_43_68 ( BL68, BLN68, WL43);
sram_cell_6t_3 inst_cell_43_67 ( BL67, BLN67, WL43);
sram_cell_6t_3 inst_cell_43_66 ( BL66, BLN66, WL43);
sram_cell_6t_3 inst_cell_43_65 ( BL65, BLN65, WL43);
sram_cell_6t_3 inst_cell_43_64 ( BL64, BLN64, WL43);
sram_cell_6t_3 inst_cell_43_63 ( BL63, BLN63, WL43);
sram_cell_6t_3 inst_cell_43_62 ( BL62, BLN62, WL43);
sram_cell_6t_3 inst_cell_43_61 ( BL61, BLN61, WL43);
sram_cell_6t_3 inst_cell_43_60 ( BL60, BLN60, WL43);
sram_cell_6t_3 inst_cell_43_59 ( BL59, BLN59, WL43);
sram_cell_6t_3 inst_cell_43_58 ( BL58, BLN58, WL43);
sram_cell_6t_3 inst_cell_43_57 ( BL57, BLN57, WL43);
sram_cell_6t_3 inst_cell_43_56 ( BL56, BLN56, WL43);
sram_cell_6t_3 inst_cell_43_55 ( BL55, BLN55, WL43);
sram_cell_6t_3 inst_cell_43_54 ( BL54, BLN54, WL43);
sram_cell_6t_3 inst_cell_43_53 ( BL53, BLN53, WL43);
sram_cell_6t_3 inst_cell_43_52 ( BL52, BLN52, WL43);
sram_cell_6t_3 inst_cell_43_51 ( BL51, BLN51, WL43);
sram_cell_6t_3 inst_cell_43_50 ( BL50, BLN50, WL43);
sram_cell_6t_3 inst_cell_43_49 ( BL49, BLN49, WL43);
sram_cell_6t_3 inst_cell_43_48 ( BL48, BLN48, WL43);
sram_cell_6t_3 inst_cell_43_47 ( BL47, BLN47, WL43);
sram_cell_6t_3 inst_cell_43_46 ( BL46, BLN46, WL43);
sram_cell_6t_3 inst_cell_43_45 ( BL45, BLN45, WL43);
sram_cell_6t_3 inst_cell_43_44 ( BL44, BLN44, WL43);
sram_cell_6t_3 inst_cell_43_43 ( BL43, BLN43, WL43);
sram_cell_6t_3 inst_cell_43_42 ( BL42, BLN42, WL43);
sram_cell_6t_3 inst_cell_43_41 ( BL41, BLN41, WL43);
sram_cell_6t_3 inst_cell_43_40 ( BL40, BLN40, WL43);
sram_cell_6t_3 inst_cell_43_39 ( BL39, BLN39, WL43);
sram_cell_6t_3 inst_cell_43_38 ( BL38, BLN38, WL43);
sram_cell_6t_3 inst_cell_43_37 ( BL37, BLN37, WL43);
sram_cell_6t_3 inst_cell_43_36 ( BL36, BLN36, WL43);
sram_cell_6t_3 inst_cell_43_35 ( BL35, BLN35, WL43);
sram_cell_6t_3 inst_cell_43_34 ( BL34, BLN34, WL43);
sram_cell_6t_3 inst_cell_43_33 ( BL33, BLN33, WL43);
sram_cell_6t_3 inst_cell_43_32 ( BL32, BLN32, WL43);
sram_cell_6t_3 inst_cell_43_31 ( BL31, BLN31, WL43);
sram_cell_6t_3 inst_cell_43_30 ( BL30, BLN30, WL43);
sram_cell_6t_3 inst_cell_43_29 ( BL29, BLN29, WL43);
sram_cell_6t_3 inst_cell_43_28 ( BL28, BLN28, WL43);
sram_cell_6t_3 inst_cell_43_27 ( BL27, BLN27, WL43);
sram_cell_6t_3 inst_cell_43_26 ( BL26, BLN26, WL43);
sram_cell_6t_3 inst_cell_43_25 ( BL25, BLN25, WL43);
sram_cell_6t_3 inst_cell_43_24 ( BL24, BLN24, WL43);
sram_cell_6t_3 inst_cell_43_23 ( BL23, BLN23, WL43);
sram_cell_6t_3 inst_cell_43_22 ( BL22, BLN22, WL43);
sram_cell_6t_3 inst_cell_43_21 ( BL21, BLN21, WL43);
sram_cell_6t_3 inst_cell_43_20 ( BL20, BLN20, WL43);
sram_cell_6t_3 inst_cell_43_19 ( BL19, BLN19, WL43);
sram_cell_6t_3 inst_cell_43_18 ( BL18, BLN18, WL43);
sram_cell_6t_3 inst_cell_43_17 ( BL17, BLN17, WL43);
sram_cell_6t_3 inst_cell_43_16 ( BL16, BLN16, WL43);
sram_cell_6t_3 inst_cell_43_15 ( BL15, BLN15, WL43);
sram_cell_6t_3 inst_cell_43_14 ( BL14, BLN14, WL43);
sram_cell_6t_3 inst_cell_43_13 ( BL13, BLN13, WL43);
sram_cell_6t_3 inst_cell_43_12 ( BL12, BLN12, WL43);
sram_cell_6t_3 inst_cell_43_11 ( BL11, BLN11, WL43);
sram_cell_6t_3 inst_cell_43_10 ( BL10, BLN10, WL43);
sram_cell_6t_3 inst_cell_43_9 ( BL9, BLN9, WL43);
sram_cell_6t_3 inst_cell_43_8 ( BL8, BLN8, WL43);
sram_cell_6t_3 inst_cell_43_7 ( BL7, BLN7, WL43);
sram_cell_6t_3 inst_cell_43_6 ( BL6, BLN6, WL43);
sram_cell_6t_3 inst_cell_43_5 ( BL5, BLN5, WL43);
sram_cell_6t_3 inst_cell_43_4 ( BL4, BLN4, WL43);
sram_cell_6t_3 inst_cell_43_3 ( BL3, BLN3, WL43);
sram_cell_6t_3 inst_cell_43_2 ( BL2, BLN2, WL43);
sram_cell_6t_3 inst_cell_43_1 ( BL1, BLN1, WL43);
sram_cell_6t_3 inst_cell_43_0 ( BL0, BLN0, WL43);
sram_cell_6t_3 inst_cell_42_127 ( BL127, BLN127, WL42);
sram_cell_6t_3 inst_cell_42_126 ( BL126, BLN126, WL42);
sram_cell_6t_3 inst_cell_42_125 ( BL125, BLN125, WL42);
sram_cell_6t_3 inst_cell_42_124 ( BL124, BLN124, WL42);
sram_cell_6t_3 inst_cell_42_123 ( BL123, BLN123, WL42);
sram_cell_6t_3 inst_cell_42_122 ( BL122, BLN122, WL42);
sram_cell_6t_3 inst_cell_42_121 ( BL121, BLN121, WL42);
sram_cell_6t_3 inst_cell_42_120 ( BL120, BLN120, WL42);
sram_cell_6t_3 inst_cell_42_119 ( BL119, BLN119, WL42);
sram_cell_6t_3 inst_cell_42_118 ( BL118, BLN118, WL42);
sram_cell_6t_3 inst_cell_42_117 ( BL117, BLN117, WL42);
sram_cell_6t_3 inst_cell_42_116 ( BL116, BLN116, WL42);
sram_cell_6t_3 inst_cell_42_115 ( BL115, BLN115, WL42);
sram_cell_6t_3 inst_cell_42_114 ( BL114, BLN114, WL42);
sram_cell_6t_3 inst_cell_42_113 ( BL113, BLN113, WL42);
sram_cell_6t_3 inst_cell_42_112 ( BL112, BLN112, WL42);
sram_cell_6t_3 inst_cell_42_111 ( BL111, BLN111, WL42);
sram_cell_6t_3 inst_cell_42_110 ( BL110, BLN110, WL42);
sram_cell_6t_3 inst_cell_42_109 ( BL109, BLN109, WL42);
sram_cell_6t_3 inst_cell_42_108 ( BL108, BLN108, WL42);
sram_cell_6t_3 inst_cell_42_107 ( BL107, BLN107, WL42);
sram_cell_6t_3 inst_cell_42_106 ( BL106, BLN106, WL42);
sram_cell_6t_3 inst_cell_42_105 ( BL105, BLN105, WL42);
sram_cell_6t_3 inst_cell_42_104 ( BL104, BLN104, WL42);
sram_cell_6t_3 inst_cell_42_103 ( BL103, BLN103, WL42);
sram_cell_6t_3 inst_cell_42_102 ( BL102, BLN102, WL42);
sram_cell_6t_3 inst_cell_42_101 ( BL101, BLN101, WL42);
sram_cell_6t_3 inst_cell_42_100 ( BL100, BLN100, WL42);
sram_cell_6t_3 inst_cell_42_99 ( BL99, BLN99, WL42);
sram_cell_6t_3 inst_cell_42_98 ( BL98, BLN98, WL42);
sram_cell_6t_3 inst_cell_42_97 ( BL97, BLN97, WL42);
sram_cell_6t_3 inst_cell_42_96 ( BL96, BLN96, WL42);
sram_cell_6t_3 inst_cell_42_95 ( BL95, BLN95, WL42);
sram_cell_6t_3 inst_cell_42_94 ( BL94, BLN94, WL42);
sram_cell_6t_3 inst_cell_42_93 ( BL93, BLN93, WL42);
sram_cell_6t_3 inst_cell_42_92 ( BL92, BLN92, WL42);
sram_cell_6t_3 inst_cell_42_91 ( BL91, BLN91, WL42);
sram_cell_6t_3 inst_cell_42_90 ( BL90, BLN90, WL42);
sram_cell_6t_3 inst_cell_42_89 ( BL89, BLN89, WL42);
sram_cell_6t_3 inst_cell_42_88 ( BL88, BLN88, WL42);
sram_cell_6t_3 inst_cell_42_87 ( BL87, BLN87, WL42);
sram_cell_6t_3 inst_cell_42_86 ( BL86, BLN86, WL42);
sram_cell_6t_3 inst_cell_42_85 ( BL85, BLN85, WL42);
sram_cell_6t_3 inst_cell_42_84 ( BL84, BLN84, WL42);
sram_cell_6t_3 inst_cell_42_83 ( BL83, BLN83, WL42);
sram_cell_6t_3 inst_cell_42_82 ( BL82, BLN82, WL42);
sram_cell_6t_3 inst_cell_42_81 ( BL81, BLN81, WL42);
sram_cell_6t_3 inst_cell_42_80 ( BL80, BLN80, WL42);
sram_cell_6t_3 inst_cell_42_79 ( BL79, BLN79, WL42);
sram_cell_6t_3 inst_cell_42_78 ( BL78, BLN78, WL42);
sram_cell_6t_3 inst_cell_42_77 ( BL77, BLN77, WL42);
sram_cell_6t_3 inst_cell_42_76 ( BL76, BLN76, WL42);
sram_cell_6t_3 inst_cell_42_75 ( BL75, BLN75, WL42);
sram_cell_6t_3 inst_cell_42_74 ( BL74, BLN74, WL42);
sram_cell_6t_3 inst_cell_42_73 ( BL73, BLN73, WL42);
sram_cell_6t_3 inst_cell_42_72 ( BL72, BLN72, WL42);
sram_cell_6t_3 inst_cell_42_71 ( BL71, BLN71, WL42);
sram_cell_6t_3 inst_cell_42_70 ( BL70, BLN70, WL42);
sram_cell_6t_3 inst_cell_42_69 ( BL69, BLN69, WL42);
sram_cell_6t_3 inst_cell_42_68 ( BL68, BLN68, WL42);
sram_cell_6t_3 inst_cell_42_67 ( BL67, BLN67, WL42);
sram_cell_6t_3 inst_cell_42_66 ( BL66, BLN66, WL42);
sram_cell_6t_3 inst_cell_42_65 ( BL65, BLN65, WL42);
sram_cell_6t_3 inst_cell_42_64 ( BL64, BLN64, WL42);
sram_cell_6t_3 inst_cell_42_63 ( BL63, BLN63, WL42);
sram_cell_6t_3 inst_cell_42_62 ( BL62, BLN62, WL42);
sram_cell_6t_3 inst_cell_42_61 ( BL61, BLN61, WL42);
sram_cell_6t_3 inst_cell_42_60 ( BL60, BLN60, WL42);
sram_cell_6t_3 inst_cell_42_59 ( BL59, BLN59, WL42);
sram_cell_6t_3 inst_cell_42_58 ( BL58, BLN58, WL42);
sram_cell_6t_3 inst_cell_42_57 ( BL57, BLN57, WL42);
sram_cell_6t_3 inst_cell_42_56 ( BL56, BLN56, WL42);
sram_cell_6t_3 inst_cell_42_55 ( BL55, BLN55, WL42);
sram_cell_6t_3 inst_cell_42_54 ( BL54, BLN54, WL42);
sram_cell_6t_3 inst_cell_42_53 ( BL53, BLN53, WL42);
sram_cell_6t_3 inst_cell_42_52 ( BL52, BLN52, WL42);
sram_cell_6t_3 inst_cell_42_51 ( BL51, BLN51, WL42);
sram_cell_6t_3 inst_cell_42_50 ( BL50, BLN50, WL42);
sram_cell_6t_3 inst_cell_42_49 ( BL49, BLN49, WL42);
sram_cell_6t_3 inst_cell_42_48 ( BL48, BLN48, WL42);
sram_cell_6t_3 inst_cell_42_47 ( BL47, BLN47, WL42);
sram_cell_6t_3 inst_cell_42_46 ( BL46, BLN46, WL42);
sram_cell_6t_3 inst_cell_42_45 ( BL45, BLN45, WL42);
sram_cell_6t_3 inst_cell_42_44 ( BL44, BLN44, WL42);
sram_cell_6t_3 inst_cell_42_43 ( BL43, BLN43, WL42);
sram_cell_6t_3 inst_cell_42_42 ( BL42, BLN42, WL42);
sram_cell_6t_3 inst_cell_42_41 ( BL41, BLN41, WL42);
sram_cell_6t_3 inst_cell_42_40 ( BL40, BLN40, WL42);
sram_cell_6t_3 inst_cell_42_39 ( BL39, BLN39, WL42);
sram_cell_6t_3 inst_cell_42_38 ( BL38, BLN38, WL42);
sram_cell_6t_3 inst_cell_42_37 ( BL37, BLN37, WL42);
sram_cell_6t_3 inst_cell_42_36 ( BL36, BLN36, WL42);
sram_cell_6t_3 inst_cell_42_35 ( BL35, BLN35, WL42);
sram_cell_6t_3 inst_cell_42_34 ( BL34, BLN34, WL42);
sram_cell_6t_3 inst_cell_42_33 ( BL33, BLN33, WL42);
sram_cell_6t_3 inst_cell_42_32 ( BL32, BLN32, WL42);
sram_cell_6t_3 inst_cell_42_31 ( BL31, BLN31, WL42);
sram_cell_6t_3 inst_cell_42_30 ( BL30, BLN30, WL42);
sram_cell_6t_3 inst_cell_42_29 ( BL29, BLN29, WL42);
sram_cell_6t_3 inst_cell_42_28 ( BL28, BLN28, WL42);
sram_cell_6t_3 inst_cell_42_27 ( BL27, BLN27, WL42);
sram_cell_6t_3 inst_cell_42_26 ( BL26, BLN26, WL42);
sram_cell_6t_3 inst_cell_42_25 ( BL25, BLN25, WL42);
sram_cell_6t_3 inst_cell_42_24 ( BL24, BLN24, WL42);
sram_cell_6t_3 inst_cell_42_23 ( BL23, BLN23, WL42);
sram_cell_6t_3 inst_cell_42_22 ( BL22, BLN22, WL42);
sram_cell_6t_3 inst_cell_42_21 ( BL21, BLN21, WL42);
sram_cell_6t_3 inst_cell_42_20 ( BL20, BLN20, WL42);
sram_cell_6t_3 inst_cell_42_19 ( BL19, BLN19, WL42);
sram_cell_6t_3 inst_cell_42_18 ( BL18, BLN18, WL42);
sram_cell_6t_3 inst_cell_42_17 ( BL17, BLN17, WL42);
sram_cell_6t_3 inst_cell_42_16 ( BL16, BLN16, WL42);
sram_cell_6t_3 inst_cell_42_15 ( BL15, BLN15, WL42);
sram_cell_6t_3 inst_cell_42_14 ( BL14, BLN14, WL42);
sram_cell_6t_3 inst_cell_42_13 ( BL13, BLN13, WL42);
sram_cell_6t_3 inst_cell_42_12 ( BL12, BLN12, WL42);
sram_cell_6t_3 inst_cell_42_11 ( BL11, BLN11, WL42);
sram_cell_6t_3 inst_cell_42_10 ( BL10, BLN10, WL42);
sram_cell_6t_3 inst_cell_42_9 ( BL9, BLN9, WL42);
sram_cell_6t_3 inst_cell_42_8 ( BL8, BLN8, WL42);
sram_cell_6t_3 inst_cell_42_7 ( BL7, BLN7, WL42);
sram_cell_6t_3 inst_cell_42_6 ( BL6, BLN6, WL42);
sram_cell_6t_3 inst_cell_42_5 ( BL5, BLN5, WL42);
sram_cell_6t_3 inst_cell_42_4 ( BL4, BLN4, WL42);
sram_cell_6t_3 inst_cell_42_3 ( BL3, BLN3, WL42);
sram_cell_6t_3 inst_cell_42_2 ( BL2, BLN2, WL42);
sram_cell_6t_3 inst_cell_42_1 ( BL1, BLN1, WL42);
sram_cell_6t_3 inst_cell_42_0 ( BL0, BLN0, WL42);
sram_cell_6t_3 inst_cell_41_127 ( BL127, BLN127, WL41);
sram_cell_6t_3 inst_cell_41_126 ( BL126, BLN126, WL41);
sram_cell_6t_3 inst_cell_41_125 ( BL125, BLN125, WL41);
sram_cell_6t_3 inst_cell_41_124 ( BL124, BLN124, WL41);
sram_cell_6t_3 inst_cell_41_123 ( BL123, BLN123, WL41);
sram_cell_6t_3 inst_cell_41_122 ( BL122, BLN122, WL41);
sram_cell_6t_3 inst_cell_41_121 ( BL121, BLN121, WL41);
sram_cell_6t_3 inst_cell_41_120 ( BL120, BLN120, WL41);
sram_cell_6t_3 inst_cell_41_119 ( BL119, BLN119, WL41);
sram_cell_6t_3 inst_cell_41_118 ( BL118, BLN118, WL41);
sram_cell_6t_3 inst_cell_41_117 ( BL117, BLN117, WL41);
sram_cell_6t_3 inst_cell_41_116 ( BL116, BLN116, WL41);
sram_cell_6t_3 inst_cell_41_115 ( BL115, BLN115, WL41);
sram_cell_6t_3 inst_cell_41_114 ( BL114, BLN114, WL41);
sram_cell_6t_3 inst_cell_41_113 ( BL113, BLN113, WL41);
sram_cell_6t_3 inst_cell_41_112 ( BL112, BLN112, WL41);
sram_cell_6t_3 inst_cell_41_111 ( BL111, BLN111, WL41);
sram_cell_6t_3 inst_cell_41_110 ( BL110, BLN110, WL41);
sram_cell_6t_3 inst_cell_41_109 ( BL109, BLN109, WL41);
sram_cell_6t_3 inst_cell_41_108 ( BL108, BLN108, WL41);
sram_cell_6t_3 inst_cell_41_107 ( BL107, BLN107, WL41);
sram_cell_6t_3 inst_cell_41_106 ( BL106, BLN106, WL41);
sram_cell_6t_3 inst_cell_41_105 ( BL105, BLN105, WL41);
sram_cell_6t_3 inst_cell_41_104 ( BL104, BLN104, WL41);
sram_cell_6t_3 inst_cell_41_103 ( BL103, BLN103, WL41);
sram_cell_6t_3 inst_cell_41_102 ( BL102, BLN102, WL41);
sram_cell_6t_3 inst_cell_41_101 ( BL101, BLN101, WL41);
sram_cell_6t_3 inst_cell_41_100 ( BL100, BLN100, WL41);
sram_cell_6t_3 inst_cell_41_99 ( BL99, BLN99, WL41);
sram_cell_6t_3 inst_cell_41_98 ( BL98, BLN98, WL41);
sram_cell_6t_3 inst_cell_41_97 ( BL97, BLN97, WL41);
sram_cell_6t_3 inst_cell_41_96 ( BL96, BLN96, WL41);
sram_cell_6t_3 inst_cell_41_95 ( BL95, BLN95, WL41);
sram_cell_6t_3 inst_cell_41_94 ( BL94, BLN94, WL41);
sram_cell_6t_3 inst_cell_41_93 ( BL93, BLN93, WL41);
sram_cell_6t_3 inst_cell_41_92 ( BL92, BLN92, WL41);
sram_cell_6t_3 inst_cell_41_91 ( BL91, BLN91, WL41);
sram_cell_6t_3 inst_cell_41_90 ( BL90, BLN90, WL41);
sram_cell_6t_3 inst_cell_41_89 ( BL89, BLN89, WL41);
sram_cell_6t_3 inst_cell_41_88 ( BL88, BLN88, WL41);
sram_cell_6t_3 inst_cell_41_87 ( BL87, BLN87, WL41);
sram_cell_6t_3 inst_cell_41_86 ( BL86, BLN86, WL41);
sram_cell_6t_3 inst_cell_41_85 ( BL85, BLN85, WL41);
sram_cell_6t_3 inst_cell_41_84 ( BL84, BLN84, WL41);
sram_cell_6t_3 inst_cell_41_83 ( BL83, BLN83, WL41);
sram_cell_6t_3 inst_cell_41_82 ( BL82, BLN82, WL41);
sram_cell_6t_3 inst_cell_41_81 ( BL81, BLN81, WL41);
sram_cell_6t_3 inst_cell_41_80 ( BL80, BLN80, WL41);
sram_cell_6t_3 inst_cell_41_79 ( BL79, BLN79, WL41);
sram_cell_6t_3 inst_cell_41_78 ( BL78, BLN78, WL41);
sram_cell_6t_3 inst_cell_41_77 ( BL77, BLN77, WL41);
sram_cell_6t_3 inst_cell_41_76 ( BL76, BLN76, WL41);
sram_cell_6t_3 inst_cell_41_75 ( BL75, BLN75, WL41);
sram_cell_6t_3 inst_cell_41_74 ( BL74, BLN74, WL41);
sram_cell_6t_3 inst_cell_41_73 ( BL73, BLN73, WL41);
sram_cell_6t_3 inst_cell_41_72 ( BL72, BLN72, WL41);
sram_cell_6t_3 inst_cell_41_71 ( BL71, BLN71, WL41);
sram_cell_6t_3 inst_cell_41_70 ( BL70, BLN70, WL41);
sram_cell_6t_3 inst_cell_41_69 ( BL69, BLN69, WL41);
sram_cell_6t_3 inst_cell_41_68 ( BL68, BLN68, WL41);
sram_cell_6t_3 inst_cell_41_67 ( BL67, BLN67, WL41);
sram_cell_6t_3 inst_cell_41_66 ( BL66, BLN66, WL41);
sram_cell_6t_3 inst_cell_41_65 ( BL65, BLN65, WL41);
sram_cell_6t_3 inst_cell_41_64 ( BL64, BLN64, WL41);
sram_cell_6t_3 inst_cell_41_63 ( BL63, BLN63, WL41);
sram_cell_6t_3 inst_cell_41_62 ( BL62, BLN62, WL41);
sram_cell_6t_3 inst_cell_41_61 ( BL61, BLN61, WL41);
sram_cell_6t_3 inst_cell_41_60 ( BL60, BLN60, WL41);
sram_cell_6t_3 inst_cell_41_59 ( BL59, BLN59, WL41);
sram_cell_6t_3 inst_cell_41_58 ( BL58, BLN58, WL41);
sram_cell_6t_3 inst_cell_41_57 ( BL57, BLN57, WL41);
sram_cell_6t_3 inst_cell_41_56 ( BL56, BLN56, WL41);
sram_cell_6t_3 inst_cell_41_55 ( BL55, BLN55, WL41);
sram_cell_6t_3 inst_cell_41_54 ( BL54, BLN54, WL41);
sram_cell_6t_3 inst_cell_41_53 ( BL53, BLN53, WL41);
sram_cell_6t_3 inst_cell_41_52 ( BL52, BLN52, WL41);
sram_cell_6t_3 inst_cell_41_51 ( BL51, BLN51, WL41);
sram_cell_6t_3 inst_cell_41_50 ( BL50, BLN50, WL41);
sram_cell_6t_3 inst_cell_41_49 ( BL49, BLN49, WL41);
sram_cell_6t_3 inst_cell_41_48 ( BL48, BLN48, WL41);
sram_cell_6t_3 inst_cell_41_47 ( BL47, BLN47, WL41);
sram_cell_6t_3 inst_cell_41_46 ( BL46, BLN46, WL41);
sram_cell_6t_3 inst_cell_41_45 ( BL45, BLN45, WL41);
sram_cell_6t_3 inst_cell_41_44 ( BL44, BLN44, WL41);
sram_cell_6t_3 inst_cell_41_43 ( BL43, BLN43, WL41);
sram_cell_6t_3 inst_cell_41_42 ( BL42, BLN42, WL41);
sram_cell_6t_3 inst_cell_41_41 ( BL41, BLN41, WL41);
sram_cell_6t_3 inst_cell_41_40 ( BL40, BLN40, WL41);
sram_cell_6t_3 inst_cell_41_39 ( BL39, BLN39, WL41);
sram_cell_6t_3 inst_cell_41_38 ( BL38, BLN38, WL41);
sram_cell_6t_3 inst_cell_41_37 ( BL37, BLN37, WL41);
sram_cell_6t_3 inst_cell_41_36 ( BL36, BLN36, WL41);
sram_cell_6t_3 inst_cell_41_35 ( BL35, BLN35, WL41);
sram_cell_6t_3 inst_cell_41_34 ( BL34, BLN34, WL41);
sram_cell_6t_3 inst_cell_41_33 ( BL33, BLN33, WL41);
sram_cell_6t_3 inst_cell_41_32 ( BL32, BLN32, WL41);
sram_cell_6t_3 inst_cell_41_31 ( BL31, BLN31, WL41);
sram_cell_6t_3 inst_cell_41_30 ( BL30, BLN30, WL41);
sram_cell_6t_3 inst_cell_41_29 ( BL29, BLN29, WL41);
sram_cell_6t_3 inst_cell_41_28 ( BL28, BLN28, WL41);
sram_cell_6t_3 inst_cell_41_27 ( BL27, BLN27, WL41);
sram_cell_6t_3 inst_cell_41_26 ( BL26, BLN26, WL41);
sram_cell_6t_3 inst_cell_41_25 ( BL25, BLN25, WL41);
sram_cell_6t_3 inst_cell_41_24 ( BL24, BLN24, WL41);
sram_cell_6t_3 inst_cell_41_23 ( BL23, BLN23, WL41);
sram_cell_6t_3 inst_cell_41_22 ( BL22, BLN22, WL41);
sram_cell_6t_3 inst_cell_41_21 ( BL21, BLN21, WL41);
sram_cell_6t_3 inst_cell_41_20 ( BL20, BLN20, WL41);
sram_cell_6t_3 inst_cell_41_19 ( BL19, BLN19, WL41);
sram_cell_6t_3 inst_cell_41_18 ( BL18, BLN18, WL41);
sram_cell_6t_3 inst_cell_41_17 ( BL17, BLN17, WL41);
sram_cell_6t_3 inst_cell_41_16 ( BL16, BLN16, WL41);
sram_cell_6t_3 inst_cell_41_15 ( BL15, BLN15, WL41);
sram_cell_6t_3 inst_cell_41_14 ( BL14, BLN14, WL41);
sram_cell_6t_3 inst_cell_41_13 ( BL13, BLN13, WL41);
sram_cell_6t_3 inst_cell_41_12 ( BL12, BLN12, WL41);
sram_cell_6t_3 inst_cell_41_11 ( BL11, BLN11, WL41);
sram_cell_6t_3 inst_cell_41_10 ( BL10, BLN10, WL41);
sram_cell_6t_3 inst_cell_41_9 ( BL9, BLN9, WL41);
sram_cell_6t_3 inst_cell_41_8 ( BL8, BLN8, WL41);
sram_cell_6t_3 inst_cell_41_7 ( BL7, BLN7, WL41);
sram_cell_6t_3 inst_cell_41_6 ( BL6, BLN6, WL41);
sram_cell_6t_3 inst_cell_41_5 ( BL5, BLN5, WL41);
sram_cell_6t_3 inst_cell_41_4 ( BL4, BLN4, WL41);
sram_cell_6t_3 inst_cell_41_3 ( BL3, BLN3, WL41);
sram_cell_6t_3 inst_cell_41_2 ( BL2, BLN2, WL41);
sram_cell_6t_3 inst_cell_41_1 ( BL1, BLN1, WL41);
sram_cell_6t_3 inst_cell_41_0 ( BL0, BLN0, WL41);
sram_cell_6t_3 inst_cell_40_127 ( BL127, BLN127, WL40);
sram_cell_6t_3 inst_cell_40_126 ( BL126, BLN126, WL40);
sram_cell_6t_3 inst_cell_40_125 ( BL125, BLN125, WL40);
sram_cell_6t_3 inst_cell_40_124 ( BL124, BLN124, WL40);
sram_cell_6t_3 inst_cell_40_123 ( BL123, BLN123, WL40);
sram_cell_6t_3 inst_cell_40_122 ( BL122, BLN122, WL40);
sram_cell_6t_3 inst_cell_40_121 ( BL121, BLN121, WL40);
sram_cell_6t_3 inst_cell_40_120 ( BL120, BLN120, WL40);
sram_cell_6t_3 inst_cell_40_119 ( BL119, BLN119, WL40);
sram_cell_6t_3 inst_cell_40_118 ( BL118, BLN118, WL40);
sram_cell_6t_3 inst_cell_40_117 ( BL117, BLN117, WL40);
sram_cell_6t_3 inst_cell_40_116 ( BL116, BLN116, WL40);
sram_cell_6t_3 inst_cell_40_115 ( BL115, BLN115, WL40);
sram_cell_6t_3 inst_cell_40_114 ( BL114, BLN114, WL40);
sram_cell_6t_3 inst_cell_40_113 ( BL113, BLN113, WL40);
sram_cell_6t_3 inst_cell_40_112 ( BL112, BLN112, WL40);
sram_cell_6t_3 inst_cell_40_111 ( BL111, BLN111, WL40);
sram_cell_6t_3 inst_cell_40_110 ( BL110, BLN110, WL40);
sram_cell_6t_3 inst_cell_40_109 ( BL109, BLN109, WL40);
sram_cell_6t_3 inst_cell_40_108 ( BL108, BLN108, WL40);
sram_cell_6t_3 inst_cell_40_107 ( BL107, BLN107, WL40);
sram_cell_6t_3 inst_cell_40_106 ( BL106, BLN106, WL40);
sram_cell_6t_3 inst_cell_40_105 ( BL105, BLN105, WL40);
sram_cell_6t_3 inst_cell_40_104 ( BL104, BLN104, WL40);
sram_cell_6t_3 inst_cell_40_103 ( BL103, BLN103, WL40);
sram_cell_6t_3 inst_cell_40_102 ( BL102, BLN102, WL40);
sram_cell_6t_3 inst_cell_40_101 ( BL101, BLN101, WL40);
sram_cell_6t_3 inst_cell_40_100 ( BL100, BLN100, WL40);
sram_cell_6t_3 inst_cell_40_99 ( BL99, BLN99, WL40);
sram_cell_6t_3 inst_cell_40_98 ( BL98, BLN98, WL40);
sram_cell_6t_3 inst_cell_40_97 ( BL97, BLN97, WL40);
sram_cell_6t_3 inst_cell_40_96 ( BL96, BLN96, WL40);
sram_cell_6t_3 inst_cell_40_95 ( BL95, BLN95, WL40);
sram_cell_6t_3 inst_cell_40_94 ( BL94, BLN94, WL40);
sram_cell_6t_3 inst_cell_40_93 ( BL93, BLN93, WL40);
sram_cell_6t_3 inst_cell_40_92 ( BL92, BLN92, WL40);
sram_cell_6t_3 inst_cell_40_91 ( BL91, BLN91, WL40);
sram_cell_6t_3 inst_cell_40_90 ( BL90, BLN90, WL40);
sram_cell_6t_3 inst_cell_40_89 ( BL89, BLN89, WL40);
sram_cell_6t_3 inst_cell_40_88 ( BL88, BLN88, WL40);
sram_cell_6t_3 inst_cell_40_87 ( BL87, BLN87, WL40);
sram_cell_6t_3 inst_cell_40_86 ( BL86, BLN86, WL40);
sram_cell_6t_3 inst_cell_40_85 ( BL85, BLN85, WL40);
sram_cell_6t_3 inst_cell_40_84 ( BL84, BLN84, WL40);
sram_cell_6t_3 inst_cell_40_83 ( BL83, BLN83, WL40);
sram_cell_6t_3 inst_cell_40_82 ( BL82, BLN82, WL40);
sram_cell_6t_3 inst_cell_40_81 ( BL81, BLN81, WL40);
sram_cell_6t_3 inst_cell_40_80 ( BL80, BLN80, WL40);
sram_cell_6t_3 inst_cell_40_79 ( BL79, BLN79, WL40);
sram_cell_6t_3 inst_cell_40_78 ( BL78, BLN78, WL40);
sram_cell_6t_3 inst_cell_40_77 ( BL77, BLN77, WL40);
sram_cell_6t_3 inst_cell_40_76 ( BL76, BLN76, WL40);
sram_cell_6t_3 inst_cell_40_75 ( BL75, BLN75, WL40);
sram_cell_6t_3 inst_cell_40_74 ( BL74, BLN74, WL40);
sram_cell_6t_3 inst_cell_40_73 ( BL73, BLN73, WL40);
sram_cell_6t_3 inst_cell_40_72 ( BL72, BLN72, WL40);
sram_cell_6t_3 inst_cell_40_71 ( BL71, BLN71, WL40);
sram_cell_6t_3 inst_cell_40_70 ( BL70, BLN70, WL40);
sram_cell_6t_3 inst_cell_40_69 ( BL69, BLN69, WL40);
sram_cell_6t_3 inst_cell_40_68 ( BL68, BLN68, WL40);
sram_cell_6t_3 inst_cell_40_67 ( BL67, BLN67, WL40);
sram_cell_6t_3 inst_cell_40_66 ( BL66, BLN66, WL40);
sram_cell_6t_3 inst_cell_40_65 ( BL65, BLN65, WL40);
sram_cell_6t_3 inst_cell_40_64 ( BL64, BLN64, WL40);
sram_cell_6t_3 inst_cell_40_63 ( BL63, BLN63, WL40);
sram_cell_6t_3 inst_cell_40_62 ( BL62, BLN62, WL40);
sram_cell_6t_3 inst_cell_40_61 ( BL61, BLN61, WL40);
sram_cell_6t_3 inst_cell_40_60 ( BL60, BLN60, WL40);
sram_cell_6t_3 inst_cell_40_59 ( BL59, BLN59, WL40);
sram_cell_6t_3 inst_cell_40_58 ( BL58, BLN58, WL40);
sram_cell_6t_3 inst_cell_40_57 ( BL57, BLN57, WL40);
sram_cell_6t_3 inst_cell_40_56 ( BL56, BLN56, WL40);
sram_cell_6t_3 inst_cell_40_55 ( BL55, BLN55, WL40);
sram_cell_6t_3 inst_cell_40_54 ( BL54, BLN54, WL40);
sram_cell_6t_3 inst_cell_40_53 ( BL53, BLN53, WL40);
sram_cell_6t_3 inst_cell_40_52 ( BL52, BLN52, WL40);
sram_cell_6t_3 inst_cell_40_51 ( BL51, BLN51, WL40);
sram_cell_6t_3 inst_cell_40_50 ( BL50, BLN50, WL40);
sram_cell_6t_3 inst_cell_40_49 ( BL49, BLN49, WL40);
sram_cell_6t_3 inst_cell_40_48 ( BL48, BLN48, WL40);
sram_cell_6t_3 inst_cell_40_47 ( BL47, BLN47, WL40);
sram_cell_6t_3 inst_cell_40_46 ( BL46, BLN46, WL40);
sram_cell_6t_3 inst_cell_40_45 ( BL45, BLN45, WL40);
sram_cell_6t_3 inst_cell_40_44 ( BL44, BLN44, WL40);
sram_cell_6t_3 inst_cell_40_43 ( BL43, BLN43, WL40);
sram_cell_6t_3 inst_cell_40_42 ( BL42, BLN42, WL40);
sram_cell_6t_3 inst_cell_40_41 ( BL41, BLN41, WL40);
sram_cell_6t_3 inst_cell_40_40 ( BL40, BLN40, WL40);
sram_cell_6t_3 inst_cell_40_39 ( BL39, BLN39, WL40);
sram_cell_6t_3 inst_cell_40_38 ( BL38, BLN38, WL40);
sram_cell_6t_3 inst_cell_40_37 ( BL37, BLN37, WL40);
sram_cell_6t_3 inst_cell_40_36 ( BL36, BLN36, WL40);
sram_cell_6t_3 inst_cell_40_35 ( BL35, BLN35, WL40);
sram_cell_6t_3 inst_cell_40_34 ( BL34, BLN34, WL40);
sram_cell_6t_3 inst_cell_40_33 ( BL33, BLN33, WL40);
sram_cell_6t_3 inst_cell_40_32 ( BL32, BLN32, WL40);
sram_cell_6t_3 inst_cell_40_31 ( BL31, BLN31, WL40);
sram_cell_6t_3 inst_cell_40_30 ( BL30, BLN30, WL40);
sram_cell_6t_3 inst_cell_40_29 ( BL29, BLN29, WL40);
sram_cell_6t_3 inst_cell_40_28 ( BL28, BLN28, WL40);
sram_cell_6t_3 inst_cell_40_27 ( BL27, BLN27, WL40);
sram_cell_6t_3 inst_cell_40_26 ( BL26, BLN26, WL40);
sram_cell_6t_3 inst_cell_40_25 ( BL25, BLN25, WL40);
sram_cell_6t_3 inst_cell_40_24 ( BL24, BLN24, WL40);
sram_cell_6t_3 inst_cell_40_23 ( BL23, BLN23, WL40);
sram_cell_6t_3 inst_cell_40_22 ( BL22, BLN22, WL40);
sram_cell_6t_3 inst_cell_40_21 ( BL21, BLN21, WL40);
sram_cell_6t_3 inst_cell_40_20 ( BL20, BLN20, WL40);
sram_cell_6t_3 inst_cell_40_19 ( BL19, BLN19, WL40);
sram_cell_6t_3 inst_cell_40_18 ( BL18, BLN18, WL40);
sram_cell_6t_3 inst_cell_40_17 ( BL17, BLN17, WL40);
sram_cell_6t_3 inst_cell_40_16 ( BL16, BLN16, WL40);
sram_cell_6t_3 inst_cell_40_15 ( BL15, BLN15, WL40);
sram_cell_6t_3 inst_cell_40_14 ( BL14, BLN14, WL40);
sram_cell_6t_3 inst_cell_40_13 ( BL13, BLN13, WL40);
sram_cell_6t_3 inst_cell_40_12 ( BL12, BLN12, WL40);
sram_cell_6t_3 inst_cell_40_11 ( BL11, BLN11, WL40);
sram_cell_6t_3 inst_cell_40_10 ( BL10, BLN10, WL40);
sram_cell_6t_3 inst_cell_40_9 ( BL9, BLN9, WL40);
sram_cell_6t_3 inst_cell_40_8 ( BL8, BLN8, WL40);
sram_cell_6t_3 inst_cell_40_7 ( BL7, BLN7, WL40);
sram_cell_6t_3 inst_cell_40_6 ( BL6, BLN6, WL40);
sram_cell_6t_3 inst_cell_40_5 ( BL5, BLN5, WL40);
sram_cell_6t_3 inst_cell_40_4 ( BL4, BLN4, WL40);
sram_cell_6t_3 inst_cell_40_3 ( BL3, BLN3, WL40);
sram_cell_6t_3 inst_cell_40_2 ( BL2, BLN2, WL40);
sram_cell_6t_3 inst_cell_40_1 ( BL1, BLN1, WL40);
sram_cell_6t_3 inst_cell_40_0 ( BL0, BLN0, WL40);
sram_cell_6t_3 inst_cell_39_127 ( BL127, BLN127, WL39);
sram_cell_6t_3 inst_cell_39_126 ( BL126, BLN126, WL39);
sram_cell_6t_3 inst_cell_39_125 ( BL125, BLN125, WL39);
sram_cell_6t_3 inst_cell_39_124 ( BL124, BLN124, WL39);
sram_cell_6t_3 inst_cell_39_123 ( BL123, BLN123, WL39);
sram_cell_6t_3 inst_cell_39_122 ( BL122, BLN122, WL39);
sram_cell_6t_3 inst_cell_39_121 ( BL121, BLN121, WL39);
sram_cell_6t_3 inst_cell_39_120 ( BL120, BLN120, WL39);
sram_cell_6t_3 inst_cell_39_119 ( BL119, BLN119, WL39);
sram_cell_6t_3 inst_cell_39_118 ( BL118, BLN118, WL39);
sram_cell_6t_3 inst_cell_39_117 ( BL117, BLN117, WL39);
sram_cell_6t_3 inst_cell_39_116 ( BL116, BLN116, WL39);
sram_cell_6t_3 inst_cell_39_115 ( BL115, BLN115, WL39);
sram_cell_6t_3 inst_cell_39_114 ( BL114, BLN114, WL39);
sram_cell_6t_3 inst_cell_39_113 ( BL113, BLN113, WL39);
sram_cell_6t_3 inst_cell_39_112 ( BL112, BLN112, WL39);
sram_cell_6t_3 inst_cell_39_111 ( BL111, BLN111, WL39);
sram_cell_6t_3 inst_cell_39_110 ( BL110, BLN110, WL39);
sram_cell_6t_3 inst_cell_39_109 ( BL109, BLN109, WL39);
sram_cell_6t_3 inst_cell_39_108 ( BL108, BLN108, WL39);
sram_cell_6t_3 inst_cell_39_107 ( BL107, BLN107, WL39);
sram_cell_6t_3 inst_cell_39_106 ( BL106, BLN106, WL39);
sram_cell_6t_3 inst_cell_39_105 ( BL105, BLN105, WL39);
sram_cell_6t_3 inst_cell_39_104 ( BL104, BLN104, WL39);
sram_cell_6t_3 inst_cell_39_103 ( BL103, BLN103, WL39);
sram_cell_6t_3 inst_cell_39_102 ( BL102, BLN102, WL39);
sram_cell_6t_3 inst_cell_39_101 ( BL101, BLN101, WL39);
sram_cell_6t_3 inst_cell_39_100 ( BL100, BLN100, WL39);
sram_cell_6t_3 inst_cell_39_99 ( BL99, BLN99, WL39);
sram_cell_6t_3 inst_cell_39_98 ( BL98, BLN98, WL39);
sram_cell_6t_3 inst_cell_39_97 ( BL97, BLN97, WL39);
sram_cell_6t_3 inst_cell_39_96 ( BL96, BLN96, WL39);
sram_cell_6t_3 inst_cell_39_95 ( BL95, BLN95, WL39);
sram_cell_6t_3 inst_cell_39_94 ( BL94, BLN94, WL39);
sram_cell_6t_3 inst_cell_39_93 ( BL93, BLN93, WL39);
sram_cell_6t_3 inst_cell_39_92 ( BL92, BLN92, WL39);
sram_cell_6t_3 inst_cell_39_91 ( BL91, BLN91, WL39);
sram_cell_6t_3 inst_cell_39_90 ( BL90, BLN90, WL39);
sram_cell_6t_3 inst_cell_39_89 ( BL89, BLN89, WL39);
sram_cell_6t_3 inst_cell_39_88 ( BL88, BLN88, WL39);
sram_cell_6t_3 inst_cell_39_87 ( BL87, BLN87, WL39);
sram_cell_6t_3 inst_cell_39_86 ( BL86, BLN86, WL39);
sram_cell_6t_3 inst_cell_39_85 ( BL85, BLN85, WL39);
sram_cell_6t_3 inst_cell_39_84 ( BL84, BLN84, WL39);
sram_cell_6t_3 inst_cell_39_83 ( BL83, BLN83, WL39);
sram_cell_6t_3 inst_cell_39_82 ( BL82, BLN82, WL39);
sram_cell_6t_3 inst_cell_39_81 ( BL81, BLN81, WL39);
sram_cell_6t_3 inst_cell_39_80 ( BL80, BLN80, WL39);
sram_cell_6t_3 inst_cell_39_79 ( BL79, BLN79, WL39);
sram_cell_6t_3 inst_cell_39_78 ( BL78, BLN78, WL39);
sram_cell_6t_3 inst_cell_39_77 ( BL77, BLN77, WL39);
sram_cell_6t_3 inst_cell_39_76 ( BL76, BLN76, WL39);
sram_cell_6t_3 inst_cell_39_75 ( BL75, BLN75, WL39);
sram_cell_6t_3 inst_cell_39_74 ( BL74, BLN74, WL39);
sram_cell_6t_3 inst_cell_39_73 ( BL73, BLN73, WL39);
sram_cell_6t_3 inst_cell_39_72 ( BL72, BLN72, WL39);
sram_cell_6t_3 inst_cell_39_71 ( BL71, BLN71, WL39);
sram_cell_6t_3 inst_cell_39_70 ( BL70, BLN70, WL39);
sram_cell_6t_3 inst_cell_39_69 ( BL69, BLN69, WL39);
sram_cell_6t_3 inst_cell_39_68 ( BL68, BLN68, WL39);
sram_cell_6t_3 inst_cell_39_67 ( BL67, BLN67, WL39);
sram_cell_6t_3 inst_cell_39_66 ( BL66, BLN66, WL39);
sram_cell_6t_3 inst_cell_39_65 ( BL65, BLN65, WL39);
sram_cell_6t_3 inst_cell_39_64 ( BL64, BLN64, WL39);
sram_cell_6t_3 inst_cell_39_63 ( BL63, BLN63, WL39);
sram_cell_6t_3 inst_cell_39_62 ( BL62, BLN62, WL39);
sram_cell_6t_3 inst_cell_39_61 ( BL61, BLN61, WL39);
sram_cell_6t_3 inst_cell_39_60 ( BL60, BLN60, WL39);
sram_cell_6t_3 inst_cell_39_59 ( BL59, BLN59, WL39);
sram_cell_6t_3 inst_cell_39_58 ( BL58, BLN58, WL39);
sram_cell_6t_3 inst_cell_39_57 ( BL57, BLN57, WL39);
sram_cell_6t_3 inst_cell_39_56 ( BL56, BLN56, WL39);
sram_cell_6t_3 inst_cell_39_55 ( BL55, BLN55, WL39);
sram_cell_6t_3 inst_cell_39_54 ( BL54, BLN54, WL39);
sram_cell_6t_3 inst_cell_39_53 ( BL53, BLN53, WL39);
sram_cell_6t_3 inst_cell_39_52 ( BL52, BLN52, WL39);
sram_cell_6t_3 inst_cell_39_51 ( BL51, BLN51, WL39);
sram_cell_6t_3 inst_cell_39_50 ( BL50, BLN50, WL39);
sram_cell_6t_3 inst_cell_39_49 ( BL49, BLN49, WL39);
sram_cell_6t_3 inst_cell_39_48 ( BL48, BLN48, WL39);
sram_cell_6t_3 inst_cell_39_47 ( BL47, BLN47, WL39);
sram_cell_6t_3 inst_cell_39_46 ( BL46, BLN46, WL39);
sram_cell_6t_3 inst_cell_39_45 ( BL45, BLN45, WL39);
sram_cell_6t_3 inst_cell_39_44 ( BL44, BLN44, WL39);
sram_cell_6t_3 inst_cell_39_43 ( BL43, BLN43, WL39);
sram_cell_6t_3 inst_cell_39_42 ( BL42, BLN42, WL39);
sram_cell_6t_3 inst_cell_39_41 ( BL41, BLN41, WL39);
sram_cell_6t_3 inst_cell_39_40 ( BL40, BLN40, WL39);
sram_cell_6t_3 inst_cell_39_39 ( BL39, BLN39, WL39);
sram_cell_6t_3 inst_cell_39_38 ( BL38, BLN38, WL39);
sram_cell_6t_3 inst_cell_39_37 ( BL37, BLN37, WL39);
sram_cell_6t_3 inst_cell_39_36 ( BL36, BLN36, WL39);
sram_cell_6t_3 inst_cell_39_35 ( BL35, BLN35, WL39);
sram_cell_6t_3 inst_cell_39_34 ( BL34, BLN34, WL39);
sram_cell_6t_3 inst_cell_39_33 ( BL33, BLN33, WL39);
sram_cell_6t_3 inst_cell_39_32 ( BL32, BLN32, WL39);
sram_cell_6t_3 inst_cell_39_31 ( BL31, BLN31, WL39);
sram_cell_6t_3 inst_cell_39_30 ( BL30, BLN30, WL39);
sram_cell_6t_3 inst_cell_39_29 ( BL29, BLN29, WL39);
sram_cell_6t_3 inst_cell_39_28 ( BL28, BLN28, WL39);
sram_cell_6t_3 inst_cell_39_27 ( BL27, BLN27, WL39);
sram_cell_6t_3 inst_cell_39_26 ( BL26, BLN26, WL39);
sram_cell_6t_3 inst_cell_39_25 ( BL25, BLN25, WL39);
sram_cell_6t_3 inst_cell_39_24 ( BL24, BLN24, WL39);
sram_cell_6t_3 inst_cell_39_23 ( BL23, BLN23, WL39);
sram_cell_6t_3 inst_cell_39_22 ( BL22, BLN22, WL39);
sram_cell_6t_3 inst_cell_39_21 ( BL21, BLN21, WL39);
sram_cell_6t_3 inst_cell_39_20 ( BL20, BLN20, WL39);
sram_cell_6t_3 inst_cell_39_19 ( BL19, BLN19, WL39);
sram_cell_6t_3 inst_cell_39_18 ( BL18, BLN18, WL39);
sram_cell_6t_3 inst_cell_39_17 ( BL17, BLN17, WL39);
sram_cell_6t_3 inst_cell_39_16 ( BL16, BLN16, WL39);
sram_cell_6t_3 inst_cell_39_15 ( BL15, BLN15, WL39);
sram_cell_6t_3 inst_cell_39_14 ( BL14, BLN14, WL39);
sram_cell_6t_3 inst_cell_39_13 ( BL13, BLN13, WL39);
sram_cell_6t_3 inst_cell_39_12 ( BL12, BLN12, WL39);
sram_cell_6t_3 inst_cell_39_11 ( BL11, BLN11, WL39);
sram_cell_6t_3 inst_cell_39_10 ( BL10, BLN10, WL39);
sram_cell_6t_3 inst_cell_39_9 ( BL9, BLN9, WL39);
sram_cell_6t_3 inst_cell_39_8 ( BL8, BLN8, WL39);
sram_cell_6t_3 inst_cell_39_7 ( BL7, BLN7, WL39);
sram_cell_6t_3 inst_cell_39_6 ( BL6, BLN6, WL39);
sram_cell_6t_3 inst_cell_39_5 ( BL5, BLN5, WL39);
sram_cell_6t_3 inst_cell_39_4 ( BL4, BLN4, WL39);
sram_cell_6t_3 inst_cell_39_3 ( BL3, BLN3, WL39);
sram_cell_6t_3 inst_cell_39_2 ( BL2, BLN2, WL39);
sram_cell_6t_3 inst_cell_39_1 ( BL1, BLN1, WL39);
sram_cell_6t_3 inst_cell_39_0 ( BL0, BLN0, WL39);
sram_cell_6t_3 inst_cell_38_127 ( BL127, BLN127, WL38);
sram_cell_6t_3 inst_cell_38_126 ( BL126, BLN126, WL38);
sram_cell_6t_3 inst_cell_38_125 ( BL125, BLN125, WL38);
sram_cell_6t_3 inst_cell_38_124 ( BL124, BLN124, WL38);
sram_cell_6t_3 inst_cell_38_123 ( BL123, BLN123, WL38);
sram_cell_6t_3 inst_cell_38_122 ( BL122, BLN122, WL38);
sram_cell_6t_3 inst_cell_38_121 ( BL121, BLN121, WL38);
sram_cell_6t_3 inst_cell_38_120 ( BL120, BLN120, WL38);
sram_cell_6t_3 inst_cell_38_119 ( BL119, BLN119, WL38);
sram_cell_6t_3 inst_cell_38_118 ( BL118, BLN118, WL38);
sram_cell_6t_3 inst_cell_38_117 ( BL117, BLN117, WL38);
sram_cell_6t_3 inst_cell_38_116 ( BL116, BLN116, WL38);
sram_cell_6t_3 inst_cell_38_115 ( BL115, BLN115, WL38);
sram_cell_6t_3 inst_cell_38_114 ( BL114, BLN114, WL38);
sram_cell_6t_3 inst_cell_38_113 ( BL113, BLN113, WL38);
sram_cell_6t_3 inst_cell_38_112 ( BL112, BLN112, WL38);
sram_cell_6t_3 inst_cell_38_111 ( BL111, BLN111, WL38);
sram_cell_6t_3 inst_cell_38_110 ( BL110, BLN110, WL38);
sram_cell_6t_3 inst_cell_38_109 ( BL109, BLN109, WL38);
sram_cell_6t_3 inst_cell_38_108 ( BL108, BLN108, WL38);
sram_cell_6t_3 inst_cell_38_107 ( BL107, BLN107, WL38);
sram_cell_6t_3 inst_cell_38_106 ( BL106, BLN106, WL38);
sram_cell_6t_3 inst_cell_38_105 ( BL105, BLN105, WL38);
sram_cell_6t_3 inst_cell_38_104 ( BL104, BLN104, WL38);
sram_cell_6t_3 inst_cell_38_103 ( BL103, BLN103, WL38);
sram_cell_6t_3 inst_cell_38_102 ( BL102, BLN102, WL38);
sram_cell_6t_3 inst_cell_38_101 ( BL101, BLN101, WL38);
sram_cell_6t_3 inst_cell_38_100 ( BL100, BLN100, WL38);
sram_cell_6t_3 inst_cell_38_99 ( BL99, BLN99, WL38);
sram_cell_6t_3 inst_cell_38_98 ( BL98, BLN98, WL38);
sram_cell_6t_3 inst_cell_38_97 ( BL97, BLN97, WL38);
sram_cell_6t_3 inst_cell_38_96 ( BL96, BLN96, WL38);
sram_cell_6t_3 inst_cell_38_95 ( BL95, BLN95, WL38);
sram_cell_6t_3 inst_cell_38_94 ( BL94, BLN94, WL38);
sram_cell_6t_3 inst_cell_38_93 ( BL93, BLN93, WL38);
sram_cell_6t_3 inst_cell_38_92 ( BL92, BLN92, WL38);
sram_cell_6t_3 inst_cell_38_91 ( BL91, BLN91, WL38);
sram_cell_6t_3 inst_cell_38_90 ( BL90, BLN90, WL38);
sram_cell_6t_3 inst_cell_38_89 ( BL89, BLN89, WL38);
sram_cell_6t_3 inst_cell_38_88 ( BL88, BLN88, WL38);
sram_cell_6t_3 inst_cell_38_87 ( BL87, BLN87, WL38);
sram_cell_6t_3 inst_cell_38_86 ( BL86, BLN86, WL38);
sram_cell_6t_3 inst_cell_38_85 ( BL85, BLN85, WL38);
sram_cell_6t_3 inst_cell_38_84 ( BL84, BLN84, WL38);
sram_cell_6t_3 inst_cell_38_83 ( BL83, BLN83, WL38);
sram_cell_6t_3 inst_cell_38_82 ( BL82, BLN82, WL38);
sram_cell_6t_3 inst_cell_38_81 ( BL81, BLN81, WL38);
sram_cell_6t_3 inst_cell_38_80 ( BL80, BLN80, WL38);
sram_cell_6t_3 inst_cell_38_79 ( BL79, BLN79, WL38);
sram_cell_6t_3 inst_cell_38_78 ( BL78, BLN78, WL38);
sram_cell_6t_3 inst_cell_38_77 ( BL77, BLN77, WL38);
sram_cell_6t_3 inst_cell_38_76 ( BL76, BLN76, WL38);
sram_cell_6t_3 inst_cell_38_75 ( BL75, BLN75, WL38);
sram_cell_6t_3 inst_cell_38_74 ( BL74, BLN74, WL38);
sram_cell_6t_3 inst_cell_38_73 ( BL73, BLN73, WL38);
sram_cell_6t_3 inst_cell_38_72 ( BL72, BLN72, WL38);
sram_cell_6t_3 inst_cell_38_71 ( BL71, BLN71, WL38);
sram_cell_6t_3 inst_cell_38_70 ( BL70, BLN70, WL38);
sram_cell_6t_3 inst_cell_38_69 ( BL69, BLN69, WL38);
sram_cell_6t_3 inst_cell_38_68 ( BL68, BLN68, WL38);
sram_cell_6t_3 inst_cell_38_67 ( BL67, BLN67, WL38);
sram_cell_6t_3 inst_cell_38_66 ( BL66, BLN66, WL38);
sram_cell_6t_3 inst_cell_38_65 ( BL65, BLN65, WL38);
sram_cell_6t_3 inst_cell_38_64 ( BL64, BLN64, WL38);
sram_cell_6t_3 inst_cell_38_63 ( BL63, BLN63, WL38);
sram_cell_6t_3 inst_cell_38_62 ( BL62, BLN62, WL38);
sram_cell_6t_3 inst_cell_38_61 ( BL61, BLN61, WL38);
sram_cell_6t_3 inst_cell_38_60 ( BL60, BLN60, WL38);
sram_cell_6t_3 inst_cell_38_59 ( BL59, BLN59, WL38);
sram_cell_6t_3 inst_cell_38_58 ( BL58, BLN58, WL38);
sram_cell_6t_3 inst_cell_38_57 ( BL57, BLN57, WL38);
sram_cell_6t_3 inst_cell_38_56 ( BL56, BLN56, WL38);
sram_cell_6t_3 inst_cell_38_55 ( BL55, BLN55, WL38);
sram_cell_6t_3 inst_cell_38_54 ( BL54, BLN54, WL38);
sram_cell_6t_3 inst_cell_38_53 ( BL53, BLN53, WL38);
sram_cell_6t_3 inst_cell_38_52 ( BL52, BLN52, WL38);
sram_cell_6t_3 inst_cell_38_51 ( BL51, BLN51, WL38);
sram_cell_6t_3 inst_cell_38_50 ( BL50, BLN50, WL38);
sram_cell_6t_3 inst_cell_38_49 ( BL49, BLN49, WL38);
sram_cell_6t_3 inst_cell_38_48 ( BL48, BLN48, WL38);
sram_cell_6t_3 inst_cell_38_47 ( BL47, BLN47, WL38);
sram_cell_6t_3 inst_cell_38_46 ( BL46, BLN46, WL38);
sram_cell_6t_3 inst_cell_38_45 ( BL45, BLN45, WL38);
sram_cell_6t_3 inst_cell_38_44 ( BL44, BLN44, WL38);
sram_cell_6t_3 inst_cell_38_43 ( BL43, BLN43, WL38);
sram_cell_6t_3 inst_cell_38_42 ( BL42, BLN42, WL38);
sram_cell_6t_3 inst_cell_38_41 ( BL41, BLN41, WL38);
sram_cell_6t_3 inst_cell_38_40 ( BL40, BLN40, WL38);
sram_cell_6t_3 inst_cell_38_39 ( BL39, BLN39, WL38);
sram_cell_6t_3 inst_cell_38_38 ( BL38, BLN38, WL38);
sram_cell_6t_3 inst_cell_38_37 ( BL37, BLN37, WL38);
sram_cell_6t_3 inst_cell_38_36 ( BL36, BLN36, WL38);
sram_cell_6t_3 inst_cell_38_35 ( BL35, BLN35, WL38);
sram_cell_6t_3 inst_cell_38_34 ( BL34, BLN34, WL38);
sram_cell_6t_3 inst_cell_38_33 ( BL33, BLN33, WL38);
sram_cell_6t_3 inst_cell_38_32 ( BL32, BLN32, WL38);
sram_cell_6t_3 inst_cell_38_31 ( BL31, BLN31, WL38);
sram_cell_6t_3 inst_cell_38_30 ( BL30, BLN30, WL38);
sram_cell_6t_3 inst_cell_38_29 ( BL29, BLN29, WL38);
sram_cell_6t_3 inst_cell_38_28 ( BL28, BLN28, WL38);
sram_cell_6t_3 inst_cell_38_27 ( BL27, BLN27, WL38);
sram_cell_6t_3 inst_cell_38_26 ( BL26, BLN26, WL38);
sram_cell_6t_3 inst_cell_38_25 ( BL25, BLN25, WL38);
sram_cell_6t_3 inst_cell_38_24 ( BL24, BLN24, WL38);
sram_cell_6t_3 inst_cell_38_23 ( BL23, BLN23, WL38);
sram_cell_6t_3 inst_cell_38_22 ( BL22, BLN22, WL38);
sram_cell_6t_3 inst_cell_38_21 ( BL21, BLN21, WL38);
sram_cell_6t_3 inst_cell_38_20 ( BL20, BLN20, WL38);
sram_cell_6t_3 inst_cell_38_19 ( BL19, BLN19, WL38);
sram_cell_6t_3 inst_cell_38_18 ( BL18, BLN18, WL38);
sram_cell_6t_3 inst_cell_38_17 ( BL17, BLN17, WL38);
sram_cell_6t_3 inst_cell_38_16 ( BL16, BLN16, WL38);
sram_cell_6t_3 inst_cell_38_15 ( BL15, BLN15, WL38);
sram_cell_6t_3 inst_cell_38_14 ( BL14, BLN14, WL38);
sram_cell_6t_3 inst_cell_38_13 ( BL13, BLN13, WL38);
sram_cell_6t_3 inst_cell_38_12 ( BL12, BLN12, WL38);
sram_cell_6t_3 inst_cell_38_11 ( BL11, BLN11, WL38);
sram_cell_6t_3 inst_cell_38_10 ( BL10, BLN10, WL38);
sram_cell_6t_3 inst_cell_38_9 ( BL9, BLN9, WL38);
sram_cell_6t_3 inst_cell_38_8 ( BL8, BLN8, WL38);
sram_cell_6t_3 inst_cell_38_7 ( BL7, BLN7, WL38);
sram_cell_6t_3 inst_cell_38_6 ( BL6, BLN6, WL38);
sram_cell_6t_3 inst_cell_38_5 ( BL5, BLN5, WL38);
sram_cell_6t_3 inst_cell_38_4 ( BL4, BLN4, WL38);
sram_cell_6t_3 inst_cell_38_3 ( BL3, BLN3, WL38);
sram_cell_6t_3 inst_cell_38_2 ( BL2, BLN2, WL38);
sram_cell_6t_3 inst_cell_38_1 ( BL1, BLN1, WL38);
sram_cell_6t_3 inst_cell_38_0 ( BL0, BLN0, WL38);
sram_cell_6t_3 inst_cell_37_127 ( BL127, BLN127, WL37);
sram_cell_6t_3 inst_cell_37_126 ( BL126, BLN126, WL37);
sram_cell_6t_3 inst_cell_37_125 ( BL125, BLN125, WL37);
sram_cell_6t_3 inst_cell_37_124 ( BL124, BLN124, WL37);
sram_cell_6t_3 inst_cell_37_123 ( BL123, BLN123, WL37);
sram_cell_6t_3 inst_cell_37_122 ( BL122, BLN122, WL37);
sram_cell_6t_3 inst_cell_37_121 ( BL121, BLN121, WL37);
sram_cell_6t_3 inst_cell_37_120 ( BL120, BLN120, WL37);
sram_cell_6t_3 inst_cell_37_119 ( BL119, BLN119, WL37);
sram_cell_6t_3 inst_cell_37_118 ( BL118, BLN118, WL37);
sram_cell_6t_3 inst_cell_37_117 ( BL117, BLN117, WL37);
sram_cell_6t_3 inst_cell_37_116 ( BL116, BLN116, WL37);
sram_cell_6t_3 inst_cell_37_115 ( BL115, BLN115, WL37);
sram_cell_6t_3 inst_cell_37_114 ( BL114, BLN114, WL37);
sram_cell_6t_3 inst_cell_37_113 ( BL113, BLN113, WL37);
sram_cell_6t_3 inst_cell_37_112 ( BL112, BLN112, WL37);
sram_cell_6t_3 inst_cell_37_111 ( BL111, BLN111, WL37);
sram_cell_6t_3 inst_cell_37_110 ( BL110, BLN110, WL37);
sram_cell_6t_3 inst_cell_37_109 ( BL109, BLN109, WL37);
sram_cell_6t_3 inst_cell_37_108 ( BL108, BLN108, WL37);
sram_cell_6t_3 inst_cell_37_107 ( BL107, BLN107, WL37);
sram_cell_6t_3 inst_cell_37_106 ( BL106, BLN106, WL37);
sram_cell_6t_3 inst_cell_37_105 ( BL105, BLN105, WL37);
sram_cell_6t_3 inst_cell_37_104 ( BL104, BLN104, WL37);
sram_cell_6t_3 inst_cell_37_103 ( BL103, BLN103, WL37);
sram_cell_6t_3 inst_cell_37_102 ( BL102, BLN102, WL37);
sram_cell_6t_3 inst_cell_37_101 ( BL101, BLN101, WL37);
sram_cell_6t_3 inst_cell_37_100 ( BL100, BLN100, WL37);
sram_cell_6t_3 inst_cell_37_99 ( BL99, BLN99, WL37);
sram_cell_6t_3 inst_cell_37_98 ( BL98, BLN98, WL37);
sram_cell_6t_3 inst_cell_37_97 ( BL97, BLN97, WL37);
sram_cell_6t_3 inst_cell_37_96 ( BL96, BLN96, WL37);
sram_cell_6t_3 inst_cell_37_95 ( BL95, BLN95, WL37);
sram_cell_6t_3 inst_cell_37_94 ( BL94, BLN94, WL37);
sram_cell_6t_3 inst_cell_37_93 ( BL93, BLN93, WL37);
sram_cell_6t_3 inst_cell_37_92 ( BL92, BLN92, WL37);
sram_cell_6t_3 inst_cell_37_91 ( BL91, BLN91, WL37);
sram_cell_6t_3 inst_cell_37_90 ( BL90, BLN90, WL37);
sram_cell_6t_3 inst_cell_37_89 ( BL89, BLN89, WL37);
sram_cell_6t_3 inst_cell_37_88 ( BL88, BLN88, WL37);
sram_cell_6t_3 inst_cell_37_87 ( BL87, BLN87, WL37);
sram_cell_6t_3 inst_cell_37_86 ( BL86, BLN86, WL37);
sram_cell_6t_3 inst_cell_37_85 ( BL85, BLN85, WL37);
sram_cell_6t_3 inst_cell_37_84 ( BL84, BLN84, WL37);
sram_cell_6t_3 inst_cell_37_83 ( BL83, BLN83, WL37);
sram_cell_6t_3 inst_cell_37_82 ( BL82, BLN82, WL37);
sram_cell_6t_3 inst_cell_37_81 ( BL81, BLN81, WL37);
sram_cell_6t_3 inst_cell_37_80 ( BL80, BLN80, WL37);
sram_cell_6t_3 inst_cell_37_79 ( BL79, BLN79, WL37);
sram_cell_6t_3 inst_cell_37_78 ( BL78, BLN78, WL37);
sram_cell_6t_3 inst_cell_37_77 ( BL77, BLN77, WL37);
sram_cell_6t_3 inst_cell_37_76 ( BL76, BLN76, WL37);
sram_cell_6t_3 inst_cell_37_75 ( BL75, BLN75, WL37);
sram_cell_6t_3 inst_cell_37_74 ( BL74, BLN74, WL37);
sram_cell_6t_3 inst_cell_37_73 ( BL73, BLN73, WL37);
sram_cell_6t_3 inst_cell_37_72 ( BL72, BLN72, WL37);
sram_cell_6t_3 inst_cell_37_71 ( BL71, BLN71, WL37);
sram_cell_6t_3 inst_cell_37_70 ( BL70, BLN70, WL37);
sram_cell_6t_3 inst_cell_37_69 ( BL69, BLN69, WL37);
sram_cell_6t_3 inst_cell_37_68 ( BL68, BLN68, WL37);
sram_cell_6t_3 inst_cell_37_67 ( BL67, BLN67, WL37);
sram_cell_6t_3 inst_cell_37_66 ( BL66, BLN66, WL37);
sram_cell_6t_3 inst_cell_37_65 ( BL65, BLN65, WL37);
sram_cell_6t_3 inst_cell_37_64 ( BL64, BLN64, WL37);
sram_cell_6t_3 inst_cell_37_63 ( BL63, BLN63, WL37);
sram_cell_6t_3 inst_cell_37_62 ( BL62, BLN62, WL37);
sram_cell_6t_3 inst_cell_37_61 ( BL61, BLN61, WL37);
sram_cell_6t_3 inst_cell_37_60 ( BL60, BLN60, WL37);
sram_cell_6t_3 inst_cell_37_59 ( BL59, BLN59, WL37);
sram_cell_6t_3 inst_cell_37_58 ( BL58, BLN58, WL37);
sram_cell_6t_3 inst_cell_37_57 ( BL57, BLN57, WL37);
sram_cell_6t_3 inst_cell_37_56 ( BL56, BLN56, WL37);
sram_cell_6t_3 inst_cell_37_55 ( BL55, BLN55, WL37);
sram_cell_6t_3 inst_cell_37_54 ( BL54, BLN54, WL37);
sram_cell_6t_3 inst_cell_37_53 ( BL53, BLN53, WL37);
sram_cell_6t_3 inst_cell_37_52 ( BL52, BLN52, WL37);
sram_cell_6t_3 inst_cell_37_51 ( BL51, BLN51, WL37);
sram_cell_6t_3 inst_cell_37_50 ( BL50, BLN50, WL37);
sram_cell_6t_3 inst_cell_37_49 ( BL49, BLN49, WL37);
sram_cell_6t_3 inst_cell_37_48 ( BL48, BLN48, WL37);
sram_cell_6t_3 inst_cell_37_47 ( BL47, BLN47, WL37);
sram_cell_6t_3 inst_cell_37_46 ( BL46, BLN46, WL37);
sram_cell_6t_3 inst_cell_37_45 ( BL45, BLN45, WL37);
sram_cell_6t_3 inst_cell_37_44 ( BL44, BLN44, WL37);
sram_cell_6t_3 inst_cell_37_43 ( BL43, BLN43, WL37);
sram_cell_6t_3 inst_cell_37_42 ( BL42, BLN42, WL37);
sram_cell_6t_3 inst_cell_37_41 ( BL41, BLN41, WL37);
sram_cell_6t_3 inst_cell_37_40 ( BL40, BLN40, WL37);
sram_cell_6t_3 inst_cell_37_39 ( BL39, BLN39, WL37);
sram_cell_6t_3 inst_cell_37_38 ( BL38, BLN38, WL37);
sram_cell_6t_3 inst_cell_37_37 ( BL37, BLN37, WL37);
sram_cell_6t_3 inst_cell_37_36 ( BL36, BLN36, WL37);
sram_cell_6t_3 inst_cell_37_35 ( BL35, BLN35, WL37);
sram_cell_6t_3 inst_cell_37_34 ( BL34, BLN34, WL37);
sram_cell_6t_3 inst_cell_37_33 ( BL33, BLN33, WL37);
sram_cell_6t_3 inst_cell_37_32 ( BL32, BLN32, WL37);
sram_cell_6t_3 inst_cell_37_31 ( BL31, BLN31, WL37);
sram_cell_6t_3 inst_cell_37_30 ( BL30, BLN30, WL37);
sram_cell_6t_3 inst_cell_37_29 ( BL29, BLN29, WL37);
sram_cell_6t_3 inst_cell_37_28 ( BL28, BLN28, WL37);
sram_cell_6t_3 inst_cell_37_27 ( BL27, BLN27, WL37);
sram_cell_6t_3 inst_cell_37_26 ( BL26, BLN26, WL37);
sram_cell_6t_3 inst_cell_37_25 ( BL25, BLN25, WL37);
sram_cell_6t_3 inst_cell_37_24 ( BL24, BLN24, WL37);
sram_cell_6t_3 inst_cell_37_23 ( BL23, BLN23, WL37);
sram_cell_6t_3 inst_cell_37_22 ( BL22, BLN22, WL37);
sram_cell_6t_3 inst_cell_37_21 ( BL21, BLN21, WL37);
sram_cell_6t_3 inst_cell_37_20 ( BL20, BLN20, WL37);
sram_cell_6t_3 inst_cell_37_19 ( BL19, BLN19, WL37);
sram_cell_6t_3 inst_cell_37_18 ( BL18, BLN18, WL37);
sram_cell_6t_3 inst_cell_37_17 ( BL17, BLN17, WL37);
sram_cell_6t_3 inst_cell_37_16 ( BL16, BLN16, WL37);
sram_cell_6t_3 inst_cell_37_15 ( BL15, BLN15, WL37);
sram_cell_6t_3 inst_cell_37_14 ( BL14, BLN14, WL37);
sram_cell_6t_3 inst_cell_37_13 ( BL13, BLN13, WL37);
sram_cell_6t_3 inst_cell_37_12 ( BL12, BLN12, WL37);
sram_cell_6t_3 inst_cell_37_11 ( BL11, BLN11, WL37);
sram_cell_6t_3 inst_cell_37_10 ( BL10, BLN10, WL37);
sram_cell_6t_3 inst_cell_37_9 ( BL9, BLN9, WL37);
sram_cell_6t_3 inst_cell_37_8 ( BL8, BLN8, WL37);
sram_cell_6t_3 inst_cell_37_7 ( BL7, BLN7, WL37);
sram_cell_6t_3 inst_cell_37_6 ( BL6, BLN6, WL37);
sram_cell_6t_3 inst_cell_37_5 ( BL5, BLN5, WL37);
sram_cell_6t_3 inst_cell_37_4 ( BL4, BLN4, WL37);
sram_cell_6t_3 inst_cell_37_3 ( BL3, BLN3, WL37);
sram_cell_6t_3 inst_cell_37_2 ( BL2, BLN2, WL37);
sram_cell_6t_3 inst_cell_37_1 ( BL1, BLN1, WL37);
sram_cell_6t_3 inst_cell_37_0 ( BL0, BLN0, WL37);
sram_cell_6t_3 inst_cell_36_127 ( BL127, BLN127, WL36);
sram_cell_6t_3 inst_cell_36_126 ( BL126, BLN126, WL36);
sram_cell_6t_3 inst_cell_36_125 ( BL125, BLN125, WL36);
sram_cell_6t_3 inst_cell_36_124 ( BL124, BLN124, WL36);
sram_cell_6t_3 inst_cell_36_123 ( BL123, BLN123, WL36);
sram_cell_6t_3 inst_cell_36_122 ( BL122, BLN122, WL36);
sram_cell_6t_3 inst_cell_36_121 ( BL121, BLN121, WL36);
sram_cell_6t_3 inst_cell_36_120 ( BL120, BLN120, WL36);
sram_cell_6t_3 inst_cell_36_119 ( BL119, BLN119, WL36);
sram_cell_6t_3 inst_cell_36_118 ( BL118, BLN118, WL36);
sram_cell_6t_3 inst_cell_36_117 ( BL117, BLN117, WL36);
sram_cell_6t_3 inst_cell_36_116 ( BL116, BLN116, WL36);
sram_cell_6t_3 inst_cell_36_115 ( BL115, BLN115, WL36);
sram_cell_6t_3 inst_cell_36_114 ( BL114, BLN114, WL36);
sram_cell_6t_3 inst_cell_36_113 ( BL113, BLN113, WL36);
sram_cell_6t_3 inst_cell_36_112 ( BL112, BLN112, WL36);
sram_cell_6t_3 inst_cell_36_111 ( BL111, BLN111, WL36);
sram_cell_6t_3 inst_cell_36_110 ( BL110, BLN110, WL36);
sram_cell_6t_3 inst_cell_36_109 ( BL109, BLN109, WL36);
sram_cell_6t_3 inst_cell_36_108 ( BL108, BLN108, WL36);
sram_cell_6t_3 inst_cell_36_107 ( BL107, BLN107, WL36);
sram_cell_6t_3 inst_cell_36_106 ( BL106, BLN106, WL36);
sram_cell_6t_3 inst_cell_36_105 ( BL105, BLN105, WL36);
sram_cell_6t_3 inst_cell_36_104 ( BL104, BLN104, WL36);
sram_cell_6t_3 inst_cell_36_103 ( BL103, BLN103, WL36);
sram_cell_6t_3 inst_cell_36_102 ( BL102, BLN102, WL36);
sram_cell_6t_3 inst_cell_36_101 ( BL101, BLN101, WL36);
sram_cell_6t_3 inst_cell_36_100 ( BL100, BLN100, WL36);
sram_cell_6t_3 inst_cell_36_99 ( BL99, BLN99, WL36);
sram_cell_6t_3 inst_cell_36_98 ( BL98, BLN98, WL36);
sram_cell_6t_3 inst_cell_36_97 ( BL97, BLN97, WL36);
sram_cell_6t_3 inst_cell_36_96 ( BL96, BLN96, WL36);
sram_cell_6t_3 inst_cell_36_95 ( BL95, BLN95, WL36);
sram_cell_6t_3 inst_cell_36_94 ( BL94, BLN94, WL36);
sram_cell_6t_3 inst_cell_36_93 ( BL93, BLN93, WL36);
sram_cell_6t_3 inst_cell_36_92 ( BL92, BLN92, WL36);
sram_cell_6t_3 inst_cell_36_91 ( BL91, BLN91, WL36);
sram_cell_6t_3 inst_cell_36_90 ( BL90, BLN90, WL36);
sram_cell_6t_3 inst_cell_36_89 ( BL89, BLN89, WL36);
sram_cell_6t_3 inst_cell_36_88 ( BL88, BLN88, WL36);
sram_cell_6t_3 inst_cell_36_87 ( BL87, BLN87, WL36);
sram_cell_6t_3 inst_cell_36_86 ( BL86, BLN86, WL36);
sram_cell_6t_3 inst_cell_36_85 ( BL85, BLN85, WL36);
sram_cell_6t_3 inst_cell_36_84 ( BL84, BLN84, WL36);
sram_cell_6t_3 inst_cell_36_83 ( BL83, BLN83, WL36);
sram_cell_6t_3 inst_cell_36_82 ( BL82, BLN82, WL36);
sram_cell_6t_3 inst_cell_36_81 ( BL81, BLN81, WL36);
sram_cell_6t_3 inst_cell_36_80 ( BL80, BLN80, WL36);
sram_cell_6t_3 inst_cell_36_79 ( BL79, BLN79, WL36);
sram_cell_6t_3 inst_cell_36_78 ( BL78, BLN78, WL36);
sram_cell_6t_3 inst_cell_36_77 ( BL77, BLN77, WL36);
sram_cell_6t_3 inst_cell_36_76 ( BL76, BLN76, WL36);
sram_cell_6t_3 inst_cell_36_75 ( BL75, BLN75, WL36);
sram_cell_6t_3 inst_cell_36_74 ( BL74, BLN74, WL36);
sram_cell_6t_3 inst_cell_36_73 ( BL73, BLN73, WL36);
sram_cell_6t_3 inst_cell_36_72 ( BL72, BLN72, WL36);
sram_cell_6t_3 inst_cell_36_71 ( BL71, BLN71, WL36);
sram_cell_6t_3 inst_cell_36_70 ( BL70, BLN70, WL36);
sram_cell_6t_3 inst_cell_36_69 ( BL69, BLN69, WL36);
sram_cell_6t_3 inst_cell_36_68 ( BL68, BLN68, WL36);
sram_cell_6t_3 inst_cell_36_67 ( BL67, BLN67, WL36);
sram_cell_6t_3 inst_cell_36_66 ( BL66, BLN66, WL36);
sram_cell_6t_3 inst_cell_36_65 ( BL65, BLN65, WL36);
sram_cell_6t_3 inst_cell_36_64 ( BL64, BLN64, WL36);
sram_cell_6t_3 inst_cell_36_63 ( BL63, BLN63, WL36);
sram_cell_6t_3 inst_cell_36_62 ( BL62, BLN62, WL36);
sram_cell_6t_3 inst_cell_36_61 ( BL61, BLN61, WL36);
sram_cell_6t_3 inst_cell_36_60 ( BL60, BLN60, WL36);
sram_cell_6t_3 inst_cell_36_59 ( BL59, BLN59, WL36);
sram_cell_6t_3 inst_cell_36_58 ( BL58, BLN58, WL36);
sram_cell_6t_3 inst_cell_36_57 ( BL57, BLN57, WL36);
sram_cell_6t_3 inst_cell_36_56 ( BL56, BLN56, WL36);
sram_cell_6t_3 inst_cell_36_55 ( BL55, BLN55, WL36);
sram_cell_6t_3 inst_cell_36_54 ( BL54, BLN54, WL36);
sram_cell_6t_3 inst_cell_36_53 ( BL53, BLN53, WL36);
sram_cell_6t_3 inst_cell_36_52 ( BL52, BLN52, WL36);
sram_cell_6t_3 inst_cell_36_51 ( BL51, BLN51, WL36);
sram_cell_6t_3 inst_cell_36_50 ( BL50, BLN50, WL36);
sram_cell_6t_3 inst_cell_36_49 ( BL49, BLN49, WL36);
sram_cell_6t_3 inst_cell_36_48 ( BL48, BLN48, WL36);
sram_cell_6t_3 inst_cell_36_47 ( BL47, BLN47, WL36);
sram_cell_6t_3 inst_cell_36_46 ( BL46, BLN46, WL36);
sram_cell_6t_3 inst_cell_36_45 ( BL45, BLN45, WL36);
sram_cell_6t_3 inst_cell_36_44 ( BL44, BLN44, WL36);
sram_cell_6t_3 inst_cell_36_43 ( BL43, BLN43, WL36);
sram_cell_6t_3 inst_cell_36_42 ( BL42, BLN42, WL36);
sram_cell_6t_3 inst_cell_36_41 ( BL41, BLN41, WL36);
sram_cell_6t_3 inst_cell_36_40 ( BL40, BLN40, WL36);
sram_cell_6t_3 inst_cell_36_39 ( BL39, BLN39, WL36);
sram_cell_6t_3 inst_cell_36_38 ( BL38, BLN38, WL36);
sram_cell_6t_3 inst_cell_36_37 ( BL37, BLN37, WL36);
sram_cell_6t_3 inst_cell_36_36 ( BL36, BLN36, WL36);
sram_cell_6t_3 inst_cell_36_35 ( BL35, BLN35, WL36);
sram_cell_6t_3 inst_cell_36_34 ( BL34, BLN34, WL36);
sram_cell_6t_3 inst_cell_36_33 ( BL33, BLN33, WL36);
sram_cell_6t_3 inst_cell_36_32 ( BL32, BLN32, WL36);
sram_cell_6t_3 inst_cell_36_31 ( BL31, BLN31, WL36);
sram_cell_6t_3 inst_cell_36_30 ( BL30, BLN30, WL36);
sram_cell_6t_3 inst_cell_36_29 ( BL29, BLN29, WL36);
sram_cell_6t_3 inst_cell_36_28 ( BL28, BLN28, WL36);
sram_cell_6t_3 inst_cell_36_27 ( BL27, BLN27, WL36);
sram_cell_6t_3 inst_cell_36_26 ( BL26, BLN26, WL36);
sram_cell_6t_3 inst_cell_36_25 ( BL25, BLN25, WL36);
sram_cell_6t_3 inst_cell_36_24 ( BL24, BLN24, WL36);
sram_cell_6t_3 inst_cell_36_23 ( BL23, BLN23, WL36);
sram_cell_6t_3 inst_cell_36_22 ( BL22, BLN22, WL36);
sram_cell_6t_3 inst_cell_36_21 ( BL21, BLN21, WL36);
sram_cell_6t_3 inst_cell_36_20 ( BL20, BLN20, WL36);
sram_cell_6t_3 inst_cell_36_19 ( BL19, BLN19, WL36);
sram_cell_6t_3 inst_cell_36_18 ( BL18, BLN18, WL36);
sram_cell_6t_3 inst_cell_36_17 ( BL17, BLN17, WL36);
sram_cell_6t_3 inst_cell_36_16 ( BL16, BLN16, WL36);
sram_cell_6t_3 inst_cell_36_15 ( BL15, BLN15, WL36);
sram_cell_6t_3 inst_cell_36_14 ( BL14, BLN14, WL36);
sram_cell_6t_3 inst_cell_36_13 ( BL13, BLN13, WL36);
sram_cell_6t_3 inst_cell_36_12 ( BL12, BLN12, WL36);
sram_cell_6t_3 inst_cell_36_11 ( BL11, BLN11, WL36);
sram_cell_6t_3 inst_cell_36_10 ( BL10, BLN10, WL36);
sram_cell_6t_3 inst_cell_36_9 ( BL9, BLN9, WL36);
sram_cell_6t_3 inst_cell_36_8 ( BL8, BLN8, WL36);
sram_cell_6t_3 inst_cell_36_7 ( BL7, BLN7, WL36);
sram_cell_6t_3 inst_cell_36_6 ( BL6, BLN6, WL36);
sram_cell_6t_3 inst_cell_36_5 ( BL5, BLN5, WL36);
sram_cell_6t_3 inst_cell_36_4 ( BL4, BLN4, WL36);
sram_cell_6t_3 inst_cell_36_3 ( BL3, BLN3, WL36);
sram_cell_6t_3 inst_cell_36_2 ( BL2, BLN2, WL36);
sram_cell_6t_3 inst_cell_36_1 ( BL1, BLN1, WL36);
sram_cell_6t_3 inst_cell_36_0 ( BL0, BLN0, WL36);
sram_cell_6t_3 inst_cell_35_127 ( BL127, BLN127, WL35);
sram_cell_6t_3 inst_cell_35_126 ( BL126, BLN126, WL35);
sram_cell_6t_3 inst_cell_35_125 ( BL125, BLN125, WL35);
sram_cell_6t_3 inst_cell_35_124 ( BL124, BLN124, WL35);
sram_cell_6t_3 inst_cell_35_123 ( BL123, BLN123, WL35);
sram_cell_6t_3 inst_cell_35_122 ( BL122, BLN122, WL35);
sram_cell_6t_3 inst_cell_35_121 ( BL121, BLN121, WL35);
sram_cell_6t_3 inst_cell_35_120 ( BL120, BLN120, WL35);
sram_cell_6t_3 inst_cell_35_119 ( BL119, BLN119, WL35);
sram_cell_6t_3 inst_cell_35_118 ( BL118, BLN118, WL35);
sram_cell_6t_3 inst_cell_35_117 ( BL117, BLN117, WL35);
sram_cell_6t_3 inst_cell_35_116 ( BL116, BLN116, WL35);
sram_cell_6t_3 inst_cell_35_115 ( BL115, BLN115, WL35);
sram_cell_6t_3 inst_cell_35_114 ( BL114, BLN114, WL35);
sram_cell_6t_3 inst_cell_35_113 ( BL113, BLN113, WL35);
sram_cell_6t_3 inst_cell_35_112 ( BL112, BLN112, WL35);
sram_cell_6t_3 inst_cell_35_111 ( BL111, BLN111, WL35);
sram_cell_6t_3 inst_cell_35_110 ( BL110, BLN110, WL35);
sram_cell_6t_3 inst_cell_35_109 ( BL109, BLN109, WL35);
sram_cell_6t_3 inst_cell_35_108 ( BL108, BLN108, WL35);
sram_cell_6t_3 inst_cell_35_107 ( BL107, BLN107, WL35);
sram_cell_6t_3 inst_cell_35_106 ( BL106, BLN106, WL35);
sram_cell_6t_3 inst_cell_35_105 ( BL105, BLN105, WL35);
sram_cell_6t_3 inst_cell_35_104 ( BL104, BLN104, WL35);
sram_cell_6t_3 inst_cell_35_103 ( BL103, BLN103, WL35);
sram_cell_6t_3 inst_cell_35_102 ( BL102, BLN102, WL35);
sram_cell_6t_3 inst_cell_35_101 ( BL101, BLN101, WL35);
sram_cell_6t_3 inst_cell_35_100 ( BL100, BLN100, WL35);
sram_cell_6t_3 inst_cell_35_99 ( BL99, BLN99, WL35);
sram_cell_6t_3 inst_cell_35_98 ( BL98, BLN98, WL35);
sram_cell_6t_3 inst_cell_35_97 ( BL97, BLN97, WL35);
sram_cell_6t_3 inst_cell_35_96 ( BL96, BLN96, WL35);
sram_cell_6t_3 inst_cell_35_95 ( BL95, BLN95, WL35);
sram_cell_6t_3 inst_cell_35_94 ( BL94, BLN94, WL35);
sram_cell_6t_3 inst_cell_35_93 ( BL93, BLN93, WL35);
sram_cell_6t_3 inst_cell_35_92 ( BL92, BLN92, WL35);
sram_cell_6t_3 inst_cell_35_91 ( BL91, BLN91, WL35);
sram_cell_6t_3 inst_cell_35_90 ( BL90, BLN90, WL35);
sram_cell_6t_3 inst_cell_35_89 ( BL89, BLN89, WL35);
sram_cell_6t_3 inst_cell_35_88 ( BL88, BLN88, WL35);
sram_cell_6t_3 inst_cell_35_87 ( BL87, BLN87, WL35);
sram_cell_6t_3 inst_cell_35_86 ( BL86, BLN86, WL35);
sram_cell_6t_3 inst_cell_35_85 ( BL85, BLN85, WL35);
sram_cell_6t_3 inst_cell_35_84 ( BL84, BLN84, WL35);
sram_cell_6t_3 inst_cell_35_83 ( BL83, BLN83, WL35);
sram_cell_6t_3 inst_cell_35_82 ( BL82, BLN82, WL35);
sram_cell_6t_3 inst_cell_35_81 ( BL81, BLN81, WL35);
sram_cell_6t_3 inst_cell_35_80 ( BL80, BLN80, WL35);
sram_cell_6t_3 inst_cell_35_79 ( BL79, BLN79, WL35);
sram_cell_6t_3 inst_cell_35_78 ( BL78, BLN78, WL35);
sram_cell_6t_3 inst_cell_35_77 ( BL77, BLN77, WL35);
sram_cell_6t_3 inst_cell_35_76 ( BL76, BLN76, WL35);
sram_cell_6t_3 inst_cell_35_75 ( BL75, BLN75, WL35);
sram_cell_6t_3 inst_cell_35_74 ( BL74, BLN74, WL35);
sram_cell_6t_3 inst_cell_35_73 ( BL73, BLN73, WL35);
sram_cell_6t_3 inst_cell_35_72 ( BL72, BLN72, WL35);
sram_cell_6t_3 inst_cell_35_71 ( BL71, BLN71, WL35);
sram_cell_6t_3 inst_cell_35_70 ( BL70, BLN70, WL35);
sram_cell_6t_3 inst_cell_35_69 ( BL69, BLN69, WL35);
sram_cell_6t_3 inst_cell_35_68 ( BL68, BLN68, WL35);
sram_cell_6t_3 inst_cell_35_67 ( BL67, BLN67, WL35);
sram_cell_6t_3 inst_cell_35_66 ( BL66, BLN66, WL35);
sram_cell_6t_3 inst_cell_35_65 ( BL65, BLN65, WL35);
sram_cell_6t_3 inst_cell_35_64 ( BL64, BLN64, WL35);
sram_cell_6t_3 inst_cell_35_63 ( BL63, BLN63, WL35);
sram_cell_6t_3 inst_cell_35_62 ( BL62, BLN62, WL35);
sram_cell_6t_3 inst_cell_35_61 ( BL61, BLN61, WL35);
sram_cell_6t_3 inst_cell_35_60 ( BL60, BLN60, WL35);
sram_cell_6t_3 inst_cell_35_59 ( BL59, BLN59, WL35);
sram_cell_6t_3 inst_cell_35_58 ( BL58, BLN58, WL35);
sram_cell_6t_3 inst_cell_35_57 ( BL57, BLN57, WL35);
sram_cell_6t_3 inst_cell_35_56 ( BL56, BLN56, WL35);
sram_cell_6t_3 inst_cell_35_55 ( BL55, BLN55, WL35);
sram_cell_6t_3 inst_cell_35_54 ( BL54, BLN54, WL35);
sram_cell_6t_3 inst_cell_35_53 ( BL53, BLN53, WL35);
sram_cell_6t_3 inst_cell_35_52 ( BL52, BLN52, WL35);
sram_cell_6t_3 inst_cell_35_51 ( BL51, BLN51, WL35);
sram_cell_6t_3 inst_cell_35_50 ( BL50, BLN50, WL35);
sram_cell_6t_3 inst_cell_35_49 ( BL49, BLN49, WL35);
sram_cell_6t_3 inst_cell_35_48 ( BL48, BLN48, WL35);
sram_cell_6t_3 inst_cell_35_47 ( BL47, BLN47, WL35);
sram_cell_6t_3 inst_cell_35_46 ( BL46, BLN46, WL35);
sram_cell_6t_3 inst_cell_35_45 ( BL45, BLN45, WL35);
sram_cell_6t_3 inst_cell_35_44 ( BL44, BLN44, WL35);
sram_cell_6t_3 inst_cell_35_43 ( BL43, BLN43, WL35);
sram_cell_6t_3 inst_cell_35_42 ( BL42, BLN42, WL35);
sram_cell_6t_3 inst_cell_35_41 ( BL41, BLN41, WL35);
sram_cell_6t_3 inst_cell_35_40 ( BL40, BLN40, WL35);
sram_cell_6t_3 inst_cell_35_39 ( BL39, BLN39, WL35);
sram_cell_6t_3 inst_cell_35_38 ( BL38, BLN38, WL35);
sram_cell_6t_3 inst_cell_35_37 ( BL37, BLN37, WL35);
sram_cell_6t_3 inst_cell_35_36 ( BL36, BLN36, WL35);
sram_cell_6t_3 inst_cell_35_35 ( BL35, BLN35, WL35);
sram_cell_6t_3 inst_cell_35_34 ( BL34, BLN34, WL35);
sram_cell_6t_3 inst_cell_35_33 ( BL33, BLN33, WL35);
sram_cell_6t_3 inst_cell_35_32 ( BL32, BLN32, WL35);
sram_cell_6t_3 inst_cell_35_31 ( BL31, BLN31, WL35);
sram_cell_6t_3 inst_cell_35_30 ( BL30, BLN30, WL35);
sram_cell_6t_3 inst_cell_35_29 ( BL29, BLN29, WL35);
sram_cell_6t_3 inst_cell_35_28 ( BL28, BLN28, WL35);
sram_cell_6t_3 inst_cell_35_27 ( BL27, BLN27, WL35);
sram_cell_6t_3 inst_cell_35_26 ( BL26, BLN26, WL35);
sram_cell_6t_3 inst_cell_35_25 ( BL25, BLN25, WL35);
sram_cell_6t_3 inst_cell_35_24 ( BL24, BLN24, WL35);
sram_cell_6t_3 inst_cell_35_23 ( BL23, BLN23, WL35);
sram_cell_6t_3 inst_cell_35_22 ( BL22, BLN22, WL35);
sram_cell_6t_3 inst_cell_35_21 ( BL21, BLN21, WL35);
sram_cell_6t_3 inst_cell_35_20 ( BL20, BLN20, WL35);
sram_cell_6t_3 inst_cell_35_19 ( BL19, BLN19, WL35);
sram_cell_6t_3 inst_cell_35_18 ( BL18, BLN18, WL35);
sram_cell_6t_3 inst_cell_35_17 ( BL17, BLN17, WL35);
sram_cell_6t_3 inst_cell_35_16 ( BL16, BLN16, WL35);
sram_cell_6t_3 inst_cell_35_15 ( BL15, BLN15, WL35);
sram_cell_6t_3 inst_cell_35_14 ( BL14, BLN14, WL35);
sram_cell_6t_3 inst_cell_35_13 ( BL13, BLN13, WL35);
sram_cell_6t_3 inst_cell_35_12 ( BL12, BLN12, WL35);
sram_cell_6t_3 inst_cell_35_11 ( BL11, BLN11, WL35);
sram_cell_6t_3 inst_cell_35_10 ( BL10, BLN10, WL35);
sram_cell_6t_3 inst_cell_35_9 ( BL9, BLN9, WL35);
sram_cell_6t_3 inst_cell_35_8 ( BL8, BLN8, WL35);
sram_cell_6t_3 inst_cell_35_7 ( BL7, BLN7, WL35);
sram_cell_6t_3 inst_cell_35_6 ( BL6, BLN6, WL35);
sram_cell_6t_3 inst_cell_35_5 ( BL5, BLN5, WL35);
sram_cell_6t_3 inst_cell_35_4 ( BL4, BLN4, WL35);
sram_cell_6t_3 inst_cell_35_3 ( BL3, BLN3, WL35);
sram_cell_6t_3 inst_cell_35_2 ( BL2, BLN2, WL35);
sram_cell_6t_3 inst_cell_35_1 ( BL1, BLN1, WL35);
sram_cell_6t_3 inst_cell_35_0 ( BL0, BLN0, WL35);
sram_cell_6t_3 inst_cell_34_127 ( BL127, BLN127, WL34);
sram_cell_6t_3 inst_cell_34_126 ( BL126, BLN126, WL34);
sram_cell_6t_3 inst_cell_34_125 ( BL125, BLN125, WL34);
sram_cell_6t_3 inst_cell_34_124 ( BL124, BLN124, WL34);
sram_cell_6t_3 inst_cell_34_123 ( BL123, BLN123, WL34);
sram_cell_6t_3 inst_cell_34_122 ( BL122, BLN122, WL34);
sram_cell_6t_3 inst_cell_34_121 ( BL121, BLN121, WL34);
sram_cell_6t_3 inst_cell_34_120 ( BL120, BLN120, WL34);
sram_cell_6t_3 inst_cell_34_119 ( BL119, BLN119, WL34);
sram_cell_6t_3 inst_cell_34_118 ( BL118, BLN118, WL34);
sram_cell_6t_3 inst_cell_34_117 ( BL117, BLN117, WL34);
sram_cell_6t_3 inst_cell_34_116 ( BL116, BLN116, WL34);
sram_cell_6t_3 inst_cell_34_115 ( BL115, BLN115, WL34);
sram_cell_6t_3 inst_cell_34_114 ( BL114, BLN114, WL34);
sram_cell_6t_3 inst_cell_34_113 ( BL113, BLN113, WL34);
sram_cell_6t_3 inst_cell_34_112 ( BL112, BLN112, WL34);
sram_cell_6t_3 inst_cell_34_111 ( BL111, BLN111, WL34);
sram_cell_6t_3 inst_cell_34_110 ( BL110, BLN110, WL34);
sram_cell_6t_3 inst_cell_34_109 ( BL109, BLN109, WL34);
sram_cell_6t_3 inst_cell_34_108 ( BL108, BLN108, WL34);
sram_cell_6t_3 inst_cell_34_107 ( BL107, BLN107, WL34);
sram_cell_6t_3 inst_cell_34_106 ( BL106, BLN106, WL34);
sram_cell_6t_3 inst_cell_34_105 ( BL105, BLN105, WL34);
sram_cell_6t_3 inst_cell_34_104 ( BL104, BLN104, WL34);
sram_cell_6t_3 inst_cell_34_103 ( BL103, BLN103, WL34);
sram_cell_6t_3 inst_cell_34_102 ( BL102, BLN102, WL34);
sram_cell_6t_3 inst_cell_34_101 ( BL101, BLN101, WL34);
sram_cell_6t_3 inst_cell_34_100 ( BL100, BLN100, WL34);
sram_cell_6t_3 inst_cell_34_99 ( BL99, BLN99, WL34);
sram_cell_6t_3 inst_cell_34_98 ( BL98, BLN98, WL34);
sram_cell_6t_3 inst_cell_34_97 ( BL97, BLN97, WL34);
sram_cell_6t_3 inst_cell_34_96 ( BL96, BLN96, WL34);
sram_cell_6t_3 inst_cell_34_95 ( BL95, BLN95, WL34);
sram_cell_6t_3 inst_cell_34_94 ( BL94, BLN94, WL34);
sram_cell_6t_3 inst_cell_34_93 ( BL93, BLN93, WL34);
sram_cell_6t_3 inst_cell_34_92 ( BL92, BLN92, WL34);
sram_cell_6t_3 inst_cell_34_91 ( BL91, BLN91, WL34);
sram_cell_6t_3 inst_cell_34_90 ( BL90, BLN90, WL34);
sram_cell_6t_3 inst_cell_34_89 ( BL89, BLN89, WL34);
sram_cell_6t_3 inst_cell_34_88 ( BL88, BLN88, WL34);
sram_cell_6t_3 inst_cell_34_87 ( BL87, BLN87, WL34);
sram_cell_6t_3 inst_cell_34_86 ( BL86, BLN86, WL34);
sram_cell_6t_3 inst_cell_34_85 ( BL85, BLN85, WL34);
sram_cell_6t_3 inst_cell_34_84 ( BL84, BLN84, WL34);
sram_cell_6t_3 inst_cell_34_83 ( BL83, BLN83, WL34);
sram_cell_6t_3 inst_cell_34_82 ( BL82, BLN82, WL34);
sram_cell_6t_3 inst_cell_34_81 ( BL81, BLN81, WL34);
sram_cell_6t_3 inst_cell_34_80 ( BL80, BLN80, WL34);
sram_cell_6t_3 inst_cell_34_79 ( BL79, BLN79, WL34);
sram_cell_6t_3 inst_cell_34_78 ( BL78, BLN78, WL34);
sram_cell_6t_3 inst_cell_34_77 ( BL77, BLN77, WL34);
sram_cell_6t_3 inst_cell_34_76 ( BL76, BLN76, WL34);
sram_cell_6t_3 inst_cell_34_75 ( BL75, BLN75, WL34);
sram_cell_6t_3 inst_cell_34_74 ( BL74, BLN74, WL34);
sram_cell_6t_3 inst_cell_34_73 ( BL73, BLN73, WL34);
sram_cell_6t_3 inst_cell_34_72 ( BL72, BLN72, WL34);
sram_cell_6t_3 inst_cell_34_71 ( BL71, BLN71, WL34);
sram_cell_6t_3 inst_cell_34_70 ( BL70, BLN70, WL34);
sram_cell_6t_3 inst_cell_34_69 ( BL69, BLN69, WL34);
sram_cell_6t_3 inst_cell_34_68 ( BL68, BLN68, WL34);
sram_cell_6t_3 inst_cell_34_67 ( BL67, BLN67, WL34);
sram_cell_6t_3 inst_cell_34_66 ( BL66, BLN66, WL34);
sram_cell_6t_3 inst_cell_34_65 ( BL65, BLN65, WL34);
sram_cell_6t_3 inst_cell_34_64 ( BL64, BLN64, WL34);
sram_cell_6t_3 inst_cell_34_63 ( BL63, BLN63, WL34);
sram_cell_6t_3 inst_cell_34_62 ( BL62, BLN62, WL34);
sram_cell_6t_3 inst_cell_34_61 ( BL61, BLN61, WL34);
sram_cell_6t_3 inst_cell_34_60 ( BL60, BLN60, WL34);
sram_cell_6t_3 inst_cell_34_59 ( BL59, BLN59, WL34);
sram_cell_6t_3 inst_cell_34_58 ( BL58, BLN58, WL34);
sram_cell_6t_3 inst_cell_34_57 ( BL57, BLN57, WL34);
sram_cell_6t_3 inst_cell_34_56 ( BL56, BLN56, WL34);
sram_cell_6t_3 inst_cell_34_55 ( BL55, BLN55, WL34);
sram_cell_6t_3 inst_cell_34_54 ( BL54, BLN54, WL34);
sram_cell_6t_3 inst_cell_34_53 ( BL53, BLN53, WL34);
sram_cell_6t_3 inst_cell_34_52 ( BL52, BLN52, WL34);
sram_cell_6t_3 inst_cell_34_51 ( BL51, BLN51, WL34);
sram_cell_6t_3 inst_cell_34_50 ( BL50, BLN50, WL34);
sram_cell_6t_3 inst_cell_34_49 ( BL49, BLN49, WL34);
sram_cell_6t_3 inst_cell_34_48 ( BL48, BLN48, WL34);
sram_cell_6t_3 inst_cell_34_47 ( BL47, BLN47, WL34);
sram_cell_6t_3 inst_cell_34_46 ( BL46, BLN46, WL34);
sram_cell_6t_3 inst_cell_34_45 ( BL45, BLN45, WL34);
sram_cell_6t_3 inst_cell_34_44 ( BL44, BLN44, WL34);
sram_cell_6t_3 inst_cell_34_43 ( BL43, BLN43, WL34);
sram_cell_6t_3 inst_cell_34_42 ( BL42, BLN42, WL34);
sram_cell_6t_3 inst_cell_34_41 ( BL41, BLN41, WL34);
sram_cell_6t_3 inst_cell_34_40 ( BL40, BLN40, WL34);
sram_cell_6t_3 inst_cell_34_39 ( BL39, BLN39, WL34);
sram_cell_6t_3 inst_cell_34_38 ( BL38, BLN38, WL34);
sram_cell_6t_3 inst_cell_34_37 ( BL37, BLN37, WL34);
sram_cell_6t_3 inst_cell_34_36 ( BL36, BLN36, WL34);
sram_cell_6t_3 inst_cell_34_35 ( BL35, BLN35, WL34);
sram_cell_6t_3 inst_cell_34_34 ( BL34, BLN34, WL34);
sram_cell_6t_3 inst_cell_34_33 ( BL33, BLN33, WL34);
sram_cell_6t_3 inst_cell_34_32 ( BL32, BLN32, WL34);
sram_cell_6t_3 inst_cell_34_31 ( BL31, BLN31, WL34);
sram_cell_6t_3 inst_cell_34_30 ( BL30, BLN30, WL34);
sram_cell_6t_3 inst_cell_34_29 ( BL29, BLN29, WL34);
sram_cell_6t_3 inst_cell_34_28 ( BL28, BLN28, WL34);
sram_cell_6t_3 inst_cell_34_27 ( BL27, BLN27, WL34);
sram_cell_6t_3 inst_cell_34_26 ( BL26, BLN26, WL34);
sram_cell_6t_3 inst_cell_34_25 ( BL25, BLN25, WL34);
sram_cell_6t_3 inst_cell_34_24 ( BL24, BLN24, WL34);
sram_cell_6t_3 inst_cell_34_23 ( BL23, BLN23, WL34);
sram_cell_6t_3 inst_cell_34_22 ( BL22, BLN22, WL34);
sram_cell_6t_3 inst_cell_34_21 ( BL21, BLN21, WL34);
sram_cell_6t_3 inst_cell_34_20 ( BL20, BLN20, WL34);
sram_cell_6t_3 inst_cell_34_19 ( BL19, BLN19, WL34);
sram_cell_6t_3 inst_cell_34_18 ( BL18, BLN18, WL34);
sram_cell_6t_3 inst_cell_34_17 ( BL17, BLN17, WL34);
sram_cell_6t_3 inst_cell_34_16 ( BL16, BLN16, WL34);
sram_cell_6t_3 inst_cell_34_15 ( BL15, BLN15, WL34);
sram_cell_6t_3 inst_cell_34_14 ( BL14, BLN14, WL34);
sram_cell_6t_3 inst_cell_34_13 ( BL13, BLN13, WL34);
sram_cell_6t_3 inst_cell_34_12 ( BL12, BLN12, WL34);
sram_cell_6t_3 inst_cell_34_11 ( BL11, BLN11, WL34);
sram_cell_6t_3 inst_cell_34_10 ( BL10, BLN10, WL34);
sram_cell_6t_3 inst_cell_34_9 ( BL9, BLN9, WL34);
sram_cell_6t_3 inst_cell_34_8 ( BL8, BLN8, WL34);
sram_cell_6t_3 inst_cell_34_7 ( BL7, BLN7, WL34);
sram_cell_6t_3 inst_cell_34_6 ( BL6, BLN6, WL34);
sram_cell_6t_3 inst_cell_34_5 ( BL5, BLN5, WL34);
sram_cell_6t_3 inst_cell_34_4 ( BL4, BLN4, WL34);
sram_cell_6t_3 inst_cell_34_3 ( BL3, BLN3, WL34);
sram_cell_6t_3 inst_cell_34_2 ( BL2, BLN2, WL34);
sram_cell_6t_3 inst_cell_34_1 ( BL1, BLN1, WL34);
sram_cell_6t_3 inst_cell_34_0 ( BL0, BLN0, WL34);
sram_cell_6t_3 inst_cell_33_127 ( BL127, BLN127, WL33);
sram_cell_6t_3 inst_cell_33_126 ( BL126, BLN126, WL33);
sram_cell_6t_3 inst_cell_33_125 ( BL125, BLN125, WL33);
sram_cell_6t_3 inst_cell_33_124 ( BL124, BLN124, WL33);
sram_cell_6t_3 inst_cell_33_123 ( BL123, BLN123, WL33);
sram_cell_6t_3 inst_cell_33_122 ( BL122, BLN122, WL33);
sram_cell_6t_3 inst_cell_33_121 ( BL121, BLN121, WL33);
sram_cell_6t_3 inst_cell_33_120 ( BL120, BLN120, WL33);
sram_cell_6t_3 inst_cell_33_119 ( BL119, BLN119, WL33);
sram_cell_6t_3 inst_cell_33_118 ( BL118, BLN118, WL33);
sram_cell_6t_3 inst_cell_33_117 ( BL117, BLN117, WL33);
sram_cell_6t_3 inst_cell_33_116 ( BL116, BLN116, WL33);
sram_cell_6t_3 inst_cell_33_115 ( BL115, BLN115, WL33);
sram_cell_6t_3 inst_cell_33_114 ( BL114, BLN114, WL33);
sram_cell_6t_3 inst_cell_33_113 ( BL113, BLN113, WL33);
sram_cell_6t_3 inst_cell_33_112 ( BL112, BLN112, WL33);
sram_cell_6t_3 inst_cell_33_111 ( BL111, BLN111, WL33);
sram_cell_6t_3 inst_cell_33_110 ( BL110, BLN110, WL33);
sram_cell_6t_3 inst_cell_33_109 ( BL109, BLN109, WL33);
sram_cell_6t_3 inst_cell_33_108 ( BL108, BLN108, WL33);
sram_cell_6t_3 inst_cell_33_107 ( BL107, BLN107, WL33);
sram_cell_6t_3 inst_cell_33_106 ( BL106, BLN106, WL33);
sram_cell_6t_3 inst_cell_33_105 ( BL105, BLN105, WL33);
sram_cell_6t_3 inst_cell_33_104 ( BL104, BLN104, WL33);
sram_cell_6t_3 inst_cell_33_103 ( BL103, BLN103, WL33);
sram_cell_6t_3 inst_cell_33_102 ( BL102, BLN102, WL33);
sram_cell_6t_3 inst_cell_33_101 ( BL101, BLN101, WL33);
sram_cell_6t_3 inst_cell_33_100 ( BL100, BLN100, WL33);
sram_cell_6t_3 inst_cell_33_99 ( BL99, BLN99, WL33);
sram_cell_6t_3 inst_cell_33_98 ( BL98, BLN98, WL33);
sram_cell_6t_3 inst_cell_33_97 ( BL97, BLN97, WL33);
sram_cell_6t_3 inst_cell_33_96 ( BL96, BLN96, WL33);
sram_cell_6t_3 inst_cell_33_95 ( BL95, BLN95, WL33);
sram_cell_6t_3 inst_cell_33_94 ( BL94, BLN94, WL33);
sram_cell_6t_3 inst_cell_33_93 ( BL93, BLN93, WL33);
sram_cell_6t_3 inst_cell_33_92 ( BL92, BLN92, WL33);
sram_cell_6t_3 inst_cell_33_91 ( BL91, BLN91, WL33);
sram_cell_6t_3 inst_cell_33_90 ( BL90, BLN90, WL33);
sram_cell_6t_3 inst_cell_33_89 ( BL89, BLN89, WL33);
sram_cell_6t_3 inst_cell_33_88 ( BL88, BLN88, WL33);
sram_cell_6t_3 inst_cell_33_87 ( BL87, BLN87, WL33);
sram_cell_6t_3 inst_cell_33_86 ( BL86, BLN86, WL33);
sram_cell_6t_3 inst_cell_33_85 ( BL85, BLN85, WL33);
sram_cell_6t_3 inst_cell_33_84 ( BL84, BLN84, WL33);
sram_cell_6t_3 inst_cell_33_83 ( BL83, BLN83, WL33);
sram_cell_6t_3 inst_cell_33_82 ( BL82, BLN82, WL33);
sram_cell_6t_3 inst_cell_33_81 ( BL81, BLN81, WL33);
sram_cell_6t_3 inst_cell_33_80 ( BL80, BLN80, WL33);
sram_cell_6t_3 inst_cell_33_79 ( BL79, BLN79, WL33);
sram_cell_6t_3 inst_cell_33_78 ( BL78, BLN78, WL33);
sram_cell_6t_3 inst_cell_33_77 ( BL77, BLN77, WL33);
sram_cell_6t_3 inst_cell_33_76 ( BL76, BLN76, WL33);
sram_cell_6t_3 inst_cell_33_75 ( BL75, BLN75, WL33);
sram_cell_6t_3 inst_cell_33_74 ( BL74, BLN74, WL33);
sram_cell_6t_3 inst_cell_33_73 ( BL73, BLN73, WL33);
sram_cell_6t_3 inst_cell_33_72 ( BL72, BLN72, WL33);
sram_cell_6t_3 inst_cell_33_71 ( BL71, BLN71, WL33);
sram_cell_6t_3 inst_cell_33_70 ( BL70, BLN70, WL33);
sram_cell_6t_3 inst_cell_33_69 ( BL69, BLN69, WL33);
sram_cell_6t_3 inst_cell_33_68 ( BL68, BLN68, WL33);
sram_cell_6t_3 inst_cell_33_67 ( BL67, BLN67, WL33);
sram_cell_6t_3 inst_cell_33_66 ( BL66, BLN66, WL33);
sram_cell_6t_3 inst_cell_33_65 ( BL65, BLN65, WL33);
sram_cell_6t_3 inst_cell_33_64 ( BL64, BLN64, WL33);
sram_cell_6t_3 inst_cell_33_63 ( BL63, BLN63, WL33);
sram_cell_6t_3 inst_cell_33_62 ( BL62, BLN62, WL33);
sram_cell_6t_3 inst_cell_33_61 ( BL61, BLN61, WL33);
sram_cell_6t_3 inst_cell_33_60 ( BL60, BLN60, WL33);
sram_cell_6t_3 inst_cell_33_59 ( BL59, BLN59, WL33);
sram_cell_6t_3 inst_cell_33_58 ( BL58, BLN58, WL33);
sram_cell_6t_3 inst_cell_33_57 ( BL57, BLN57, WL33);
sram_cell_6t_3 inst_cell_33_56 ( BL56, BLN56, WL33);
sram_cell_6t_3 inst_cell_33_55 ( BL55, BLN55, WL33);
sram_cell_6t_3 inst_cell_33_54 ( BL54, BLN54, WL33);
sram_cell_6t_3 inst_cell_33_53 ( BL53, BLN53, WL33);
sram_cell_6t_3 inst_cell_33_52 ( BL52, BLN52, WL33);
sram_cell_6t_3 inst_cell_33_51 ( BL51, BLN51, WL33);
sram_cell_6t_3 inst_cell_33_50 ( BL50, BLN50, WL33);
sram_cell_6t_3 inst_cell_33_49 ( BL49, BLN49, WL33);
sram_cell_6t_3 inst_cell_33_48 ( BL48, BLN48, WL33);
sram_cell_6t_3 inst_cell_33_47 ( BL47, BLN47, WL33);
sram_cell_6t_3 inst_cell_33_46 ( BL46, BLN46, WL33);
sram_cell_6t_3 inst_cell_33_45 ( BL45, BLN45, WL33);
sram_cell_6t_3 inst_cell_33_44 ( BL44, BLN44, WL33);
sram_cell_6t_3 inst_cell_33_43 ( BL43, BLN43, WL33);
sram_cell_6t_3 inst_cell_33_42 ( BL42, BLN42, WL33);
sram_cell_6t_3 inst_cell_33_41 ( BL41, BLN41, WL33);
sram_cell_6t_3 inst_cell_33_40 ( BL40, BLN40, WL33);
sram_cell_6t_3 inst_cell_33_39 ( BL39, BLN39, WL33);
sram_cell_6t_3 inst_cell_33_38 ( BL38, BLN38, WL33);
sram_cell_6t_3 inst_cell_33_37 ( BL37, BLN37, WL33);
sram_cell_6t_3 inst_cell_33_36 ( BL36, BLN36, WL33);
sram_cell_6t_3 inst_cell_33_35 ( BL35, BLN35, WL33);
sram_cell_6t_3 inst_cell_33_34 ( BL34, BLN34, WL33);
sram_cell_6t_3 inst_cell_33_33 ( BL33, BLN33, WL33);
sram_cell_6t_3 inst_cell_33_32 ( BL32, BLN32, WL33);
sram_cell_6t_3 inst_cell_33_31 ( BL31, BLN31, WL33);
sram_cell_6t_3 inst_cell_33_30 ( BL30, BLN30, WL33);
sram_cell_6t_3 inst_cell_33_29 ( BL29, BLN29, WL33);
sram_cell_6t_3 inst_cell_33_28 ( BL28, BLN28, WL33);
sram_cell_6t_3 inst_cell_33_27 ( BL27, BLN27, WL33);
sram_cell_6t_3 inst_cell_33_26 ( BL26, BLN26, WL33);
sram_cell_6t_3 inst_cell_33_25 ( BL25, BLN25, WL33);
sram_cell_6t_3 inst_cell_33_24 ( BL24, BLN24, WL33);
sram_cell_6t_3 inst_cell_33_23 ( BL23, BLN23, WL33);
sram_cell_6t_3 inst_cell_33_22 ( BL22, BLN22, WL33);
sram_cell_6t_3 inst_cell_33_21 ( BL21, BLN21, WL33);
sram_cell_6t_3 inst_cell_33_20 ( BL20, BLN20, WL33);
sram_cell_6t_3 inst_cell_33_19 ( BL19, BLN19, WL33);
sram_cell_6t_3 inst_cell_33_18 ( BL18, BLN18, WL33);
sram_cell_6t_3 inst_cell_33_17 ( BL17, BLN17, WL33);
sram_cell_6t_3 inst_cell_33_16 ( BL16, BLN16, WL33);
sram_cell_6t_3 inst_cell_33_15 ( BL15, BLN15, WL33);
sram_cell_6t_3 inst_cell_33_14 ( BL14, BLN14, WL33);
sram_cell_6t_3 inst_cell_33_13 ( BL13, BLN13, WL33);
sram_cell_6t_3 inst_cell_33_12 ( BL12, BLN12, WL33);
sram_cell_6t_3 inst_cell_33_11 ( BL11, BLN11, WL33);
sram_cell_6t_3 inst_cell_33_10 ( BL10, BLN10, WL33);
sram_cell_6t_3 inst_cell_33_9 ( BL9, BLN9, WL33);
sram_cell_6t_3 inst_cell_33_8 ( BL8, BLN8, WL33);
sram_cell_6t_3 inst_cell_33_7 ( BL7, BLN7, WL33);
sram_cell_6t_3 inst_cell_33_6 ( BL6, BLN6, WL33);
sram_cell_6t_3 inst_cell_33_5 ( BL5, BLN5, WL33);
sram_cell_6t_3 inst_cell_33_4 ( BL4, BLN4, WL33);
sram_cell_6t_3 inst_cell_33_3 ( BL3, BLN3, WL33);
sram_cell_6t_3 inst_cell_33_2 ( BL2, BLN2, WL33);
sram_cell_6t_3 inst_cell_33_1 ( BL1, BLN1, WL33);
sram_cell_6t_3 inst_cell_33_0 ( BL0, BLN0, WL33);
sram_cell_6t_3 inst_cell_32_127 ( BL127, BLN127, WL32);
sram_cell_6t_3 inst_cell_32_126 ( BL126, BLN126, WL32);
sram_cell_6t_3 inst_cell_32_125 ( BL125, BLN125, WL32);
sram_cell_6t_3 inst_cell_32_124 ( BL124, BLN124, WL32);
sram_cell_6t_3 inst_cell_32_123 ( BL123, BLN123, WL32);
sram_cell_6t_3 inst_cell_32_122 ( BL122, BLN122, WL32);
sram_cell_6t_3 inst_cell_32_121 ( BL121, BLN121, WL32);
sram_cell_6t_3 inst_cell_32_120 ( BL120, BLN120, WL32);
sram_cell_6t_3 inst_cell_32_119 ( BL119, BLN119, WL32);
sram_cell_6t_3 inst_cell_32_118 ( BL118, BLN118, WL32);
sram_cell_6t_3 inst_cell_32_117 ( BL117, BLN117, WL32);
sram_cell_6t_3 inst_cell_32_116 ( BL116, BLN116, WL32);
sram_cell_6t_3 inst_cell_32_115 ( BL115, BLN115, WL32);
sram_cell_6t_3 inst_cell_32_114 ( BL114, BLN114, WL32);
sram_cell_6t_3 inst_cell_32_113 ( BL113, BLN113, WL32);
sram_cell_6t_3 inst_cell_32_112 ( BL112, BLN112, WL32);
sram_cell_6t_3 inst_cell_32_111 ( BL111, BLN111, WL32);
sram_cell_6t_3 inst_cell_32_110 ( BL110, BLN110, WL32);
sram_cell_6t_3 inst_cell_32_109 ( BL109, BLN109, WL32);
sram_cell_6t_3 inst_cell_32_108 ( BL108, BLN108, WL32);
sram_cell_6t_3 inst_cell_32_107 ( BL107, BLN107, WL32);
sram_cell_6t_3 inst_cell_32_106 ( BL106, BLN106, WL32);
sram_cell_6t_3 inst_cell_32_105 ( BL105, BLN105, WL32);
sram_cell_6t_3 inst_cell_32_104 ( BL104, BLN104, WL32);
sram_cell_6t_3 inst_cell_32_103 ( BL103, BLN103, WL32);
sram_cell_6t_3 inst_cell_32_102 ( BL102, BLN102, WL32);
sram_cell_6t_3 inst_cell_32_101 ( BL101, BLN101, WL32);
sram_cell_6t_3 inst_cell_32_100 ( BL100, BLN100, WL32);
sram_cell_6t_3 inst_cell_32_99 ( BL99, BLN99, WL32);
sram_cell_6t_3 inst_cell_32_98 ( BL98, BLN98, WL32);
sram_cell_6t_3 inst_cell_32_97 ( BL97, BLN97, WL32);
sram_cell_6t_3 inst_cell_32_96 ( BL96, BLN96, WL32);
sram_cell_6t_3 inst_cell_32_95 ( BL95, BLN95, WL32);
sram_cell_6t_3 inst_cell_32_94 ( BL94, BLN94, WL32);
sram_cell_6t_3 inst_cell_32_93 ( BL93, BLN93, WL32);
sram_cell_6t_3 inst_cell_32_92 ( BL92, BLN92, WL32);
sram_cell_6t_3 inst_cell_32_91 ( BL91, BLN91, WL32);
sram_cell_6t_3 inst_cell_32_90 ( BL90, BLN90, WL32);
sram_cell_6t_3 inst_cell_32_89 ( BL89, BLN89, WL32);
sram_cell_6t_3 inst_cell_32_88 ( BL88, BLN88, WL32);
sram_cell_6t_3 inst_cell_32_87 ( BL87, BLN87, WL32);
sram_cell_6t_3 inst_cell_32_86 ( BL86, BLN86, WL32);
sram_cell_6t_3 inst_cell_32_85 ( BL85, BLN85, WL32);
sram_cell_6t_3 inst_cell_32_84 ( BL84, BLN84, WL32);
sram_cell_6t_3 inst_cell_32_83 ( BL83, BLN83, WL32);
sram_cell_6t_3 inst_cell_32_82 ( BL82, BLN82, WL32);
sram_cell_6t_3 inst_cell_32_81 ( BL81, BLN81, WL32);
sram_cell_6t_3 inst_cell_32_80 ( BL80, BLN80, WL32);
sram_cell_6t_3 inst_cell_32_79 ( BL79, BLN79, WL32);
sram_cell_6t_3 inst_cell_32_78 ( BL78, BLN78, WL32);
sram_cell_6t_3 inst_cell_32_77 ( BL77, BLN77, WL32);
sram_cell_6t_3 inst_cell_32_76 ( BL76, BLN76, WL32);
sram_cell_6t_3 inst_cell_32_75 ( BL75, BLN75, WL32);
sram_cell_6t_3 inst_cell_32_74 ( BL74, BLN74, WL32);
sram_cell_6t_3 inst_cell_32_73 ( BL73, BLN73, WL32);
sram_cell_6t_3 inst_cell_32_72 ( BL72, BLN72, WL32);
sram_cell_6t_3 inst_cell_32_71 ( BL71, BLN71, WL32);
sram_cell_6t_3 inst_cell_32_70 ( BL70, BLN70, WL32);
sram_cell_6t_3 inst_cell_32_69 ( BL69, BLN69, WL32);
sram_cell_6t_3 inst_cell_32_68 ( BL68, BLN68, WL32);
sram_cell_6t_3 inst_cell_32_67 ( BL67, BLN67, WL32);
sram_cell_6t_3 inst_cell_32_66 ( BL66, BLN66, WL32);
sram_cell_6t_3 inst_cell_32_65 ( BL65, BLN65, WL32);
sram_cell_6t_3 inst_cell_32_64 ( BL64, BLN64, WL32);
sram_cell_6t_3 inst_cell_32_63 ( BL63, BLN63, WL32);
sram_cell_6t_3 inst_cell_32_62 ( BL62, BLN62, WL32);
sram_cell_6t_3 inst_cell_32_61 ( BL61, BLN61, WL32);
sram_cell_6t_3 inst_cell_32_60 ( BL60, BLN60, WL32);
sram_cell_6t_3 inst_cell_32_59 ( BL59, BLN59, WL32);
sram_cell_6t_3 inst_cell_32_58 ( BL58, BLN58, WL32);
sram_cell_6t_3 inst_cell_32_57 ( BL57, BLN57, WL32);
sram_cell_6t_3 inst_cell_32_56 ( BL56, BLN56, WL32);
sram_cell_6t_3 inst_cell_32_55 ( BL55, BLN55, WL32);
sram_cell_6t_3 inst_cell_32_54 ( BL54, BLN54, WL32);
sram_cell_6t_3 inst_cell_32_53 ( BL53, BLN53, WL32);
sram_cell_6t_3 inst_cell_32_52 ( BL52, BLN52, WL32);
sram_cell_6t_3 inst_cell_32_51 ( BL51, BLN51, WL32);
sram_cell_6t_3 inst_cell_32_50 ( BL50, BLN50, WL32);
sram_cell_6t_3 inst_cell_32_49 ( BL49, BLN49, WL32);
sram_cell_6t_3 inst_cell_32_48 ( BL48, BLN48, WL32);
sram_cell_6t_3 inst_cell_32_47 ( BL47, BLN47, WL32);
sram_cell_6t_3 inst_cell_32_46 ( BL46, BLN46, WL32);
sram_cell_6t_3 inst_cell_32_45 ( BL45, BLN45, WL32);
sram_cell_6t_3 inst_cell_32_44 ( BL44, BLN44, WL32);
sram_cell_6t_3 inst_cell_32_43 ( BL43, BLN43, WL32);
sram_cell_6t_3 inst_cell_32_42 ( BL42, BLN42, WL32);
sram_cell_6t_3 inst_cell_32_41 ( BL41, BLN41, WL32);
sram_cell_6t_3 inst_cell_32_40 ( BL40, BLN40, WL32);
sram_cell_6t_3 inst_cell_32_39 ( BL39, BLN39, WL32);
sram_cell_6t_3 inst_cell_32_38 ( BL38, BLN38, WL32);
sram_cell_6t_3 inst_cell_32_37 ( BL37, BLN37, WL32);
sram_cell_6t_3 inst_cell_32_36 ( BL36, BLN36, WL32);
sram_cell_6t_3 inst_cell_32_35 ( BL35, BLN35, WL32);
sram_cell_6t_3 inst_cell_32_34 ( BL34, BLN34, WL32);
sram_cell_6t_3 inst_cell_32_33 ( BL33, BLN33, WL32);
sram_cell_6t_3 inst_cell_32_32 ( BL32, BLN32, WL32);
sram_cell_6t_3 inst_cell_32_31 ( BL31, BLN31, WL32);
sram_cell_6t_3 inst_cell_32_30 ( BL30, BLN30, WL32);
sram_cell_6t_3 inst_cell_32_29 ( BL29, BLN29, WL32);
sram_cell_6t_3 inst_cell_32_28 ( BL28, BLN28, WL32);
sram_cell_6t_3 inst_cell_32_27 ( BL27, BLN27, WL32);
sram_cell_6t_3 inst_cell_32_26 ( BL26, BLN26, WL32);
sram_cell_6t_3 inst_cell_32_25 ( BL25, BLN25, WL32);
sram_cell_6t_3 inst_cell_32_24 ( BL24, BLN24, WL32);
sram_cell_6t_3 inst_cell_32_23 ( BL23, BLN23, WL32);
sram_cell_6t_3 inst_cell_32_22 ( BL22, BLN22, WL32);
sram_cell_6t_3 inst_cell_32_21 ( BL21, BLN21, WL32);
sram_cell_6t_3 inst_cell_32_20 ( BL20, BLN20, WL32);
sram_cell_6t_3 inst_cell_32_19 ( BL19, BLN19, WL32);
sram_cell_6t_3 inst_cell_32_18 ( BL18, BLN18, WL32);
sram_cell_6t_3 inst_cell_32_17 ( BL17, BLN17, WL32);
sram_cell_6t_3 inst_cell_32_16 ( BL16, BLN16, WL32);
sram_cell_6t_3 inst_cell_32_15 ( BL15, BLN15, WL32);
sram_cell_6t_3 inst_cell_32_14 ( BL14, BLN14, WL32);
sram_cell_6t_3 inst_cell_32_13 ( BL13, BLN13, WL32);
sram_cell_6t_3 inst_cell_32_12 ( BL12, BLN12, WL32);
sram_cell_6t_3 inst_cell_32_11 ( BL11, BLN11, WL32);
sram_cell_6t_3 inst_cell_32_10 ( BL10, BLN10, WL32);
sram_cell_6t_3 inst_cell_32_9 ( BL9, BLN9, WL32);
sram_cell_6t_3 inst_cell_32_8 ( BL8, BLN8, WL32);
sram_cell_6t_3 inst_cell_32_7 ( BL7, BLN7, WL32);
sram_cell_6t_3 inst_cell_32_6 ( BL6, BLN6, WL32);
sram_cell_6t_3 inst_cell_32_5 ( BL5, BLN5, WL32);
sram_cell_6t_3 inst_cell_32_4 ( BL4, BLN4, WL32);
sram_cell_6t_3 inst_cell_32_3 ( BL3, BLN3, WL32);
sram_cell_6t_3 inst_cell_32_2 ( BL2, BLN2, WL32);
sram_cell_6t_3 inst_cell_32_1 ( BL1, BLN1, WL32);
sram_cell_6t_3 inst_cell_32_0 ( BL0, BLN0, WL32);
sram_cell_6t_3 inst_cell_31_127 ( BL127, BLN127, WL31);
sram_cell_6t_3 inst_cell_31_126 ( BL126, BLN126, WL31);
sram_cell_6t_3 inst_cell_31_125 ( BL125, BLN125, WL31);
sram_cell_6t_3 inst_cell_31_124 ( BL124, BLN124, WL31);
sram_cell_6t_3 inst_cell_31_123 ( BL123, BLN123, WL31);
sram_cell_6t_3 inst_cell_31_122 ( BL122, BLN122, WL31);
sram_cell_6t_3 inst_cell_31_121 ( BL121, BLN121, WL31);
sram_cell_6t_3 inst_cell_31_120 ( BL120, BLN120, WL31);
sram_cell_6t_3 inst_cell_31_119 ( BL119, BLN119, WL31);
sram_cell_6t_3 inst_cell_31_118 ( BL118, BLN118, WL31);
sram_cell_6t_3 inst_cell_31_117 ( BL117, BLN117, WL31);
sram_cell_6t_3 inst_cell_31_116 ( BL116, BLN116, WL31);
sram_cell_6t_3 inst_cell_31_115 ( BL115, BLN115, WL31);
sram_cell_6t_3 inst_cell_31_114 ( BL114, BLN114, WL31);
sram_cell_6t_3 inst_cell_31_113 ( BL113, BLN113, WL31);
sram_cell_6t_3 inst_cell_31_112 ( BL112, BLN112, WL31);
sram_cell_6t_3 inst_cell_31_111 ( BL111, BLN111, WL31);
sram_cell_6t_3 inst_cell_31_110 ( BL110, BLN110, WL31);
sram_cell_6t_3 inst_cell_31_109 ( BL109, BLN109, WL31);
sram_cell_6t_3 inst_cell_31_108 ( BL108, BLN108, WL31);
sram_cell_6t_3 inst_cell_31_107 ( BL107, BLN107, WL31);
sram_cell_6t_3 inst_cell_31_106 ( BL106, BLN106, WL31);
sram_cell_6t_3 inst_cell_31_105 ( BL105, BLN105, WL31);
sram_cell_6t_3 inst_cell_31_104 ( BL104, BLN104, WL31);
sram_cell_6t_3 inst_cell_31_103 ( BL103, BLN103, WL31);
sram_cell_6t_3 inst_cell_31_102 ( BL102, BLN102, WL31);
sram_cell_6t_3 inst_cell_31_101 ( BL101, BLN101, WL31);
sram_cell_6t_3 inst_cell_31_100 ( BL100, BLN100, WL31);
sram_cell_6t_3 inst_cell_31_99 ( BL99, BLN99, WL31);
sram_cell_6t_3 inst_cell_31_98 ( BL98, BLN98, WL31);
sram_cell_6t_3 inst_cell_31_97 ( BL97, BLN97, WL31);
sram_cell_6t_3 inst_cell_31_96 ( BL96, BLN96, WL31);
sram_cell_6t_3 inst_cell_31_95 ( BL95, BLN95, WL31);
sram_cell_6t_3 inst_cell_31_94 ( BL94, BLN94, WL31);
sram_cell_6t_3 inst_cell_31_93 ( BL93, BLN93, WL31);
sram_cell_6t_3 inst_cell_31_92 ( BL92, BLN92, WL31);
sram_cell_6t_3 inst_cell_31_91 ( BL91, BLN91, WL31);
sram_cell_6t_3 inst_cell_31_90 ( BL90, BLN90, WL31);
sram_cell_6t_3 inst_cell_31_89 ( BL89, BLN89, WL31);
sram_cell_6t_3 inst_cell_31_88 ( BL88, BLN88, WL31);
sram_cell_6t_3 inst_cell_31_87 ( BL87, BLN87, WL31);
sram_cell_6t_3 inst_cell_31_86 ( BL86, BLN86, WL31);
sram_cell_6t_3 inst_cell_31_85 ( BL85, BLN85, WL31);
sram_cell_6t_3 inst_cell_31_84 ( BL84, BLN84, WL31);
sram_cell_6t_3 inst_cell_31_83 ( BL83, BLN83, WL31);
sram_cell_6t_3 inst_cell_31_82 ( BL82, BLN82, WL31);
sram_cell_6t_3 inst_cell_31_81 ( BL81, BLN81, WL31);
sram_cell_6t_3 inst_cell_31_80 ( BL80, BLN80, WL31);
sram_cell_6t_3 inst_cell_31_79 ( BL79, BLN79, WL31);
sram_cell_6t_3 inst_cell_31_78 ( BL78, BLN78, WL31);
sram_cell_6t_3 inst_cell_31_77 ( BL77, BLN77, WL31);
sram_cell_6t_3 inst_cell_31_76 ( BL76, BLN76, WL31);
sram_cell_6t_3 inst_cell_31_75 ( BL75, BLN75, WL31);
sram_cell_6t_3 inst_cell_31_74 ( BL74, BLN74, WL31);
sram_cell_6t_3 inst_cell_31_73 ( BL73, BLN73, WL31);
sram_cell_6t_3 inst_cell_31_72 ( BL72, BLN72, WL31);
sram_cell_6t_3 inst_cell_31_71 ( BL71, BLN71, WL31);
sram_cell_6t_3 inst_cell_31_70 ( BL70, BLN70, WL31);
sram_cell_6t_3 inst_cell_31_69 ( BL69, BLN69, WL31);
sram_cell_6t_3 inst_cell_31_68 ( BL68, BLN68, WL31);
sram_cell_6t_3 inst_cell_31_67 ( BL67, BLN67, WL31);
sram_cell_6t_3 inst_cell_31_66 ( BL66, BLN66, WL31);
sram_cell_6t_3 inst_cell_31_65 ( BL65, BLN65, WL31);
sram_cell_6t_3 inst_cell_31_64 ( BL64, BLN64, WL31);
sram_cell_6t_3 inst_cell_31_63 ( BL63, BLN63, WL31);
sram_cell_6t_3 inst_cell_31_62 ( BL62, BLN62, WL31);
sram_cell_6t_3 inst_cell_31_61 ( BL61, BLN61, WL31);
sram_cell_6t_3 inst_cell_31_60 ( BL60, BLN60, WL31);
sram_cell_6t_3 inst_cell_31_59 ( BL59, BLN59, WL31);
sram_cell_6t_3 inst_cell_31_58 ( BL58, BLN58, WL31);
sram_cell_6t_3 inst_cell_31_57 ( BL57, BLN57, WL31);
sram_cell_6t_3 inst_cell_31_56 ( BL56, BLN56, WL31);
sram_cell_6t_3 inst_cell_31_55 ( BL55, BLN55, WL31);
sram_cell_6t_3 inst_cell_31_54 ( BL54, BLN54, WL31);
sram_cell_6t_3 inst_cell_31_53 ( BL53, BLN53, WL31);
sram_cell_6t_3 inst_cell_31_52 ( BL52, BLN52, WL31);
sram_cell_6t_3 inst_cell_31_51 ( BL51, BLN51, WL31);
sram_cell_6t_3 inst_cell_31_50 ( BL50, BLN50, WL31);
sram_cell_6t_3 inst_cell_31_49 ( BL49, BLN49, WL31);
sram_cell_6t_3 inst_cell_31_48 ( BL48, BLN48, WL31);
sram_cell_6t_3 inst_cell_31_47 ( BL47, BLN47, WL31);
sram_cell_6t_3 inst_cell_31_46 ( BL46, BLN46, WL31);
sram_cell_6t_3 inst_cell_31_45 ( BL45, BLN45, WL31);
sram_cell_6t_3 inst_cell_31_44 ( BL44, BLN44, WL31);
sram_cell_6t_3 inst_cell_31_43 ( BL43, BLN43, WL31);
sram_cell_6t_3 inst_cell_31_42 ( BL42, BLN42, WL31);
sram_cell_6t_3 inst_cell_31_41 ( BL41, BLN41, WL31);
sram_cell_6t_3 inst_cell_31_40 ( BL40, BLN40, WL31);
sram_cell_6t_3 inst_cell_31_39 ( BL39, BLN39, WL31);
sram_cell_6t_3 inst_cell_31_38 ( BL38, BLN38, WL31);
sram_cell_6t_3 inst_cell_31_37 ( BL37, BLN37, WL31);
sram_cell_6t_3 inst_cell_31_36 ( BL36, BLN36, WL31);
sram_cell_6t_3 inst_cell_31_35 ( BL35, BLN35, WL31);
sram_cell_6t_3 inst_cell_31_34 ( BL34, BLN34, WL31);
sram_cell_6t_3 inst_cell_31_33 ( BL33, BLN33, WL31);
sram_cell_6t_3 inst_cell_31_32 ( BL32, BLN32, WL31);
sram_cell_6t_3 inst_cell_31_31 ( BL31, BLN31, WL31);
sram_cell_6t_3 inst_cell_31_30 ( BL30, BLN30, WL31);
sram_cell_6t_3 inst_cell_31_29 ( BL29, BLN29, WL31);
sram_cell_6t_3 inst_cell_31_28 ( BL28, BLN28, WL31);
sram_cell_6t_3 inst_cell_31_27 ( BL27, BLN27, WL31);
sram_cell_6t_3 inst_cell_31_26 ( BL26, BLN26, WL31);
sram_cell_6t_3 inst_cell_31_25 ( BL25, BLN25, WL31);
sram_cell_6t_3 inst_cell_31_24 ( BL24, BLN24, WL31);
sram_cell_6t_3 inst_cell_31_23 ( BL23, BLN23, WL31);
sram_cell_6t_3 inst_cell_31_22 ( BL22, BLN22, WL31);
sram_cell_6t_3 inst_cell_31_21 ( BL21, BLN21, WL31);
sram_cell_6t_3 inst_cell_31_20 ( BL20, BLN20, WL31);
sram_cell_6t_3 inst_cell_31_19 ( BL19, BLN19, WL31);
sram_cell_6t_3 inst_cell_31_18 ( BL18, BLN18, WL31);
sram_cell_6t_3 inst_cell_31_17 ( BL17, BLN17, WL31);
sram_cell_6t_3 inst_cell_31_16 ( BL16, BLN16, WL31);
sram_cell_6t_3 inst_cell_31_15 ( BL15, BLN15, WL31);
sram_cell_6t_3 inst_cell_31_14 ( BL14, BLN14, WL31);
sram_cell_6t_3 inst_cell_31_13 ( BL13, BLN13, WL31);
sram_cell_6t_3 inst_cell_31_12 ( BL12, BLN12, WL31);
sram_cell_6t_3 inst_cell_31_11 ( BL11, BLN11, WL31);
sram_cell_6t_3 inst_cell_31_10 ( BL10, BLN10, WL31);
sram_cell_6t_3 inst_cell_31_9 ( BL9, BLN9, WL31);
sram_cell_6t_3 inst_cell_31_8 ( BL8, BLN8, WL31);
sram_cell_6t_3 inst_cell_31_7 ( BL7, BLN7, WL31);
sram_cell_6t_3 inst_cell_31_6 ( BL6, BLN6, WL31);
sram_cell_6t_3 inst_cell_31_5 ( BL5, BLN5, WL31);
sram_cell_6t_3 inst_cell_31_4 ( BL4, BLN4, WL31);
sram_cell_6t_3 inst_cell_31_3 ( BL3, BLN3, WL31);
sram_cell_6t_3 inst_cell_31_2 ( BL2, BLN2, WL31);
sram_cell_6t_3 inst_cell_31_1 ( BL1, BLN1, WL31);
sram_cell_6t_3 inst_cell_31_0 ( BL0, BLN0, WL31);
sram_cell_6t_3 inst_cell_30_127 ( BL127, BLN127, WL30);
sram_cell_6t_3 inst_cell_30_126 ( BL126, BLN126, WL30);
sram_cell_6t_3 inst_cell_30_125 ( BL125, BLN125, WL30);
sram_cell_6t_3 inst_cell_30_124 ( BL124, BLN124, WL30);
sram_cell_6t_3 inst_cell_30_123 ( BL123, BLN123, WL30);
sram_cell_6t_3 inst_cell_30_122 ( BL122, BLN122, WL30);
sram_cell_6t_3 inst_cell_30_121 ( BL121, BLN121, WL30);
sram_cell_6t_3 inst_cell_30_120 ( BL120, BLN120, WL30);
sram_cell_6t_3 inst_cell_30_119 ( BL119, BLN119, WL30);
sram_cell_6t_3 inst_cell_30_118 ( BL118, BLN118, WL30);
sram_cell_6t_3 inst_cell_30_117 ( BL117, BLN117, WL30);
sram_cell_6t_3 inst_cell_30_116 ( BL116, BLN116, WL30);
sram_cell_6t_3 inst_cell_30_115 ( BL115, BLN115, WL30);
sram_cell_6t_3 inst_cell_30_114 ( BL114, BLN114, WL30);
sram_cell_6t_3 inst_cell_30_113 ( BL113, BLN113, WL30);
sram_cell_6t_3 inst_cell_30_112 ( BL112, BLN112, WL30);
sram_cell_6t_3 inst_cell_30_111 ( BL111, BLN111, WL30);
sram_cell_6t_3 inst_cell_30_110 ( BL110, BLN110, WL30);
sram_cell_6t_3 inst_cell_30_109 ( BL109, BLN109, WL30);
sram_cell_6t_3 inst_cell_30_108 ( BL108, BLN108, WL30);
sram_cell_6t_3 inst_cell_30_107 ( BL107, BLN107, WL30);
sram_cell_6t_3 inst_cell_30_106 ( BL106, BLN106, WL30);
sram_cell_6t_3 inst_cell_30_105 ( BL105, BLN105, WL30);
sram_cell_6t_3 inst_cell_30_104 ( BL104, BLN104, WL30);
sram_cell_6t_3 inst_cell_30_103 ( BL103, BLN103, WL30);
sram_cell_6t_3 inst_cell_30_102 ( BL102, BLN102, WL30);
sram_cell_6t_3 inst_cell_30_101 ( BL101, BLN101, WL30);
sram_cell_6t_3 inst_cell_30_100 ( BL100, BLN100, WL30);
sram_cell_6t_3 inst_cell_30_99 ( BL99, BLN99, WL30);
sram_cell_6t_3 inst_cell_30_98 ( BL98, BLN98, WL30);
sram_cell_6t_3 inst_cell_30_97 ( BL97, BLN97, WL30);
sram_cell_6t_3 inst_cell_30_96 ( BL96, BLN96, WL30);
sram_cell_6t_3 inst_cell_30_95 ( BL95, BLN95, WL30);
sram_cell_6t_3 inst_cell_30_94 ( BL94, BLN94, WL30);
sram_cell_6t_3 inst_cell_30_93 ( BL93, BLN93, WL30);
sram_cell_6t_3 inst_cell_30_92 ( BL92, BLN92, WL30);
sram_cell_6t_3 inst_cell_30_91 ( BL91, BLN91, WL30);
sram_cell_6t_3 inst_cell_30_90 ( BL90, BLN90, WL30);
sram_cell_6t_3 inst_cell_30_89 ( BL89, BLN89, WL30);
sram_cell_6t_3 inst_cell_30_88 ( BL88, BLN88, WL30);
sram_cell_6t_3 inst_cell_30_87 ( BL87, BLN87, WL30);
sram_cell_6t_3 inst_cell_30_86 ( BL86, BLN86, WL30);
sram_cell_6t_3 inst_cell_30_85 ( BL85, BLN85, WL30);
sram_cell_6t_3 inst_cell_30_84 ( BL84, BLN84, WL30);
sram_cell_6t_3 inst_cell_30_83 ( BL83, BLN83, WL30);
sram_cell_6t_3 inst_cell_30_82 ( BL82, BLN82, WL30);
sram_cell_6t_3 inst_cell_30_81 ( BL81, BLN81, WL30);
sram_cell_6t_3 inst_cell_30_80 ( BL80, BLN80, WL30);
sram_cell_6t_3 inst_cell_30_79 ( BL79, BLN79, WL30);
sram_cell_6t_3 inst_cell_30_78 ( BL78, BLN78, WL30);
sram_cell_6t_3 inst_cell_30_77 ( BL77, BLN77, WL30);
sram_cell_6t_3 inst_cell_30_76 ( BL76, BLN76, WL30);
sram_cell_6t_3 inst_cell_30_75 ( BL75, BLN75, WL30);
sram_cell_6t_3 inst_cell_30_74 ( BL74, BLN74, WL30);
sram_cell_6t_3 inst_cell_30_73 ( BL73, BLN73, WL30);
sram_cell_6t_3 inst_cell_30_72 ( BL72, BLN72, WL30);
sram_cell_6t_3 inst_cell_30_71 ( BL71, BLN71, WL30);
sram_cell_6t_3 inst_cell_30_70 ( BL70, BLN70, WL30);
sram_cell_6t_3 inst_cell_30_69 ( BL69, BLN69, WL30);
sram_cell_6t_3 inst_cell_30_68 ( BL68, BLN68, WL30);
sram_cell_6t_3 inst_cell_30_67 ( BL67, BLN67, WL30);
sram_cell_6t_3 inst_cell_30_66 ( BL66, BLN66, WL30);
sram_cell_6t_3 inst_cell_30_65 ( BL65, BLN65, WL30);
sram_cell_6t_3 inst_cell_30_64 ( BL64, BLN64, WL30);
sram_cell_6t_3 inst_cell_30_63 ( BL63, BLN63, WL30);
sram_cell_6t_3 inst_cell_30_62 ( BL62, BLN62, WL30);
sram_cell_6t_3 inst_cell_30_61 ( BL61, BLN61, WL30);
sram_cell_6t_3 inst_cell_30_60 ( BL60, BLN60, WL30);
sram_cell_6t_3 inst_cell_30_59 ( BL59, BLN59, WL30);
sram_cell_6t_3 inst_cell_30_58 ( BL58, BLN58, WL30);
sram_cell_6t_3 inst_cell_30_57 ( BL57, BLN57, WL30);
sram_cell_6t_3 inst_cell_30_56 ( BL56, BLN56, WL30);
sram_cell_6t_3 inst_cell_30_55 ( BL55, BLN55, WL30);
sram_cell_6t_3 inst_cell_30_54 ( BL54, BLN54, WL30);
sram_cell_6t_3 inst_cell_30_53 ( BL53, BLN53, WL30);
sram_cell_6t_3 inst_cell_30_52 ( BL52, BLN52, WL30);
sram_cell_6t_3 inst_cell_30_51 ( BL51, BLN51, WL30);
sram_cell_6t_3 inst_cell_30_50 ( BL50, BLN50, WL30);
sram_cell_6t_3 inst_cell_30_49 ( BL49, BLN49, WL30);
sram_cell_6t_3 inst_cell_30_48 ( BL48, BLN48, WL30);
sram_cell_6t_3 inst_cell_30_47 ( BL47, BLN47, WL30);
sram_cell_6t_3 inst_cell_30_46 ( BL46, BLN46, WL30);
sram_cell_6t_3 inst_cell_30_45 ( BL45, BLN45, WL30);
sram_cell_6t_3 inst_cell_30_44 ( BL44, BLN44, WL30);
sram_cell_6t_3 inst_cell_30_43 ( BL43, BLN43, WL30);
sram_cell_6t_3 inst_cell_30_42 ( BL42, BLN42, WL30);
sram_cell_6t_3 inst_cell_30_41 ( BL41, BLN41, WL30);
sram_cell_6t_3 inst_cell_30_40 ( BL40, BLN40, WL30);
sram_cell_6t_3 inst_cell_30_39 ( BL39, BLN39, WL30);
sram_cell_6t_3 inst_cell_30_38 ( BL38, BLN38, WL30);
sram_cell_6t_3 inst_cell_30_37 ( BL37, BLN37, WL30);
sram_cell_6t_3 inst_cell_30_36 ( BL36, BLN36, WL30);
sram_cell_6t_3 inst_cell_30_35 ( BL35, BLN35, WL30);
sram_cell_6t_3 inst_cell_30_34 ( BL34, BLN34, WL30);
sram_cell_6t_3 inst_cell_30_33 ( BL33, BLN33, WL30);
sram_cell_6t_3 inst_cell_30_32 ( BL32, BLN32, WL30);
sram_cell_6t_3 inst_cell_30_31 ( BL31, BLN31, WL30);
sram_cell_6t_3 inst_cell_30_30 ( BL30, BLN30, WL30);
sram_cell_6t_3 inst_cell_30_29 ( BL29, BLN29, WL30);
sram_cell_6t_3 inst_cell_30_28 ( BL28, BLN28, WL30);
sram_cell_6t_3 inst_cell_30_27 ( BL27, BLN27, WL30);
sram_cell_6t_3 inst_cell_30_26 ( BL26, BLN26, WL30);
sram_cell_6t_3 inst_cell_30_25 ( BL25, BLN25, WL30);
sram_cell_6t_3 inst_cell_30_24 ( BL24, BLN24, WL30);
sram_cell_6t_3 inst_cell_30_23 ( BL23, BLN23, WL30);
sram_cell_6t_3 inst_cell_30_22 ( BL22, BLN22, WL30);
sram_cell_6t_3 inst_cell_30_21 ( BL21, BLN21, WL30);
sram_cell_6t_3 inst_cell_30_20 ( BL20, BLN20, WL30);
sram_cell_6t_3 inst_cell_30_19 ( BL19, BLN19, WL30);
sram_cell_6t_3 inst_cell_30_18 ( BL18, BLN18, WL30);
sram_cell_6t_3 inst_cell_30_17 ( BL17, BLN17, WL30);
sram_cell_6t_3 inst_cell_30_16 ( BL16, BLN16, WL30);
sram_cell_6t_3 inst_cell_30_15 ( BL15, BLN15, WL30);
sram_cell_6t_3 inst_cell_30_14 ( BL14, BLN14, WL30);
sram_cell_6t_3 inst_cell_30_13 ( BL13, BLN13, WL30);
sram_cell_6t_3 inst_cell_30_12 ( BL12, BLN12, WL30);
sram_cell_6t_3 inst_cell_30_11 ( BL11, BLN11, WL30);
sram_cell_6t_3 inst_cell_30_10 ( BL10, BLN10, WL30);
sram_cell_6t_3 inst_cell_30_9 ( BL9, BLN9, WL30);
sram_cell_6t_3 inst_cell_30_8 ( BL8, BLN8, WL30);
sram_cell_6t_3 inst_cell_30_7 ( BL7, BLN7, WL30);
sram_cell_6t_3 inst_cell_30_6 ( BL6, BLN6, WL30);
sram_cell_6t_3 inst_cell_30_5 ( BL5, BLN5, WL30);
sram_cell_6t_3 inst_cell_30_4 ( BL4, BLN4, WL30);
sram_cell_6t_3 inst_cell_30_3 ( BL3, BLN3, WL30);
sram_cell_6t_3 inst_cell_30_2 ( BL2, BLN2, WL30);
sram_cell_6t_3 inst_cell_30_1 ( BL1, BLN1, WL30);
sram_cell_6t_3 inst_cell_30_0 ( BL0, BLN0, WL30);
sram_cell_6t_3 inst_cell_29_127 ( BL127, BLN127, WL29);
sram_cell_6t_3 inst_cell_29_126 ( BL126, BLN126, WL29);
sram_cell_6t_3 inst_cell_29_125 ( BL125, BLN125, WL29);
sram_cell_6t_3 inst_cell_29_124 ( BL124, BLN124, WL29);
sram_cell_6t_3 inst_cell_29_123 ( BL123, BLN123, WL29);
sram_cell_6t_3 inst_cell_29_122 ( BL122, BLN122, WL29);
sram_cell_6t_3 inst_cell_29_121 ( BL121, BLN121, WL29);
sram_cell_6t_3 inst_cell_29_120 ( BL120, BLN120, WL29);
sram_cell_6t_3 inst_cell_29_119 ( BL119, BLN119, WL29);
sram_cell_6t_3 inst_cell_29_118 ( BL118, BLN118, WL29);
sram_cell_6t_3 inst_cell_29_117 ( BL117, BLN117, WL29);
sram_cell_6t_3 inst_cell_29_116 ( BL116, BLN116, WL29);
sram_cell_6t_3 inst_cell_29_115 ( BL115, BLN115, WL29);
sram_cell_6t_3 inst_cell_29_114 ( BL114, BLN114, WL29);
sram_cell_6t_3 inst_cell_29_113 ( BL113, BLN113, WL29);
sram_cell_6t_3 inst_cell_29_112 ( BL112, BLN112, WL29);
sram_cell_6t_3 inst_cell_29_111 ( BL111, BLN111, WL29);
sram_cell_6t_3 inst_cell_29_110 ( BL110, BLN110, WL29);
sram_cell_6t_3 inst_cell_29_109 ( BL109, BLN109, WL29);
sram_cell_6t_3 inst_cell_29_108 ( BL108, BLN108, WL29);
sram_cell_6t_3 inst_cell_29_107 ( BL107, BLN107, WL29);
sram_cell_6t_3 inst_cell_29_106 ( BL106, BLN106, WL29);
sram_cell_6t_3 inst_cell_29_105 ( BL105, BLN105, WL29);
sram_cell_6t_3 inst_cell_29_104 ( BL104, BLN104, WL29);
sram_cell_6t_3 inst_cell_29_103 ( BL103, BLN103, WL29);
sram_cell_6t_3 inst_cell_29_102 ( BL102, BLN102, WL29);
sram_cell_6t_3 inst_cell_29_101 ( BL101, BLN101, WL29);
sram_cell_6t_3 inst_cell_29_100 ( BL100, BLN100, WL29);
sram_cell_6t_3 inst_cell_29_99 ( BL99, BLN99, WL29);
sram_cell_6t_3 inst_cell_29_98 ( BL98, BLN98, WL29);
sram_cell_6t_3 inst_cell_29_97 ( BL97, BLN97, WL29);
sram_cell_6t_3 inst_cell_29_96 ( BL96, BLN96, WL29);
sram_cell_6t_3 inst_cell_29_95 ( BL95, BLN95, WL29);
sram_cell_6t_3 inst_cell_29_94 ( BL94, BLN94, WL29);
sram_cell_6t_3 inst_cell_29_93 ( BL93, BLN93, WL29);
sram_cell_6t_3 inst_cell_29_92 ( BL92, BLN92, WL29);
sram_cell_6t_3 inst_cell_29_91 ( BL91, BLN91, WL29);
sram_cell_6t_3 inst_cell_29_90 ( BL90, BLN90, WL29);
sram_cell_6t_3 inst_cell_29_89 ( BL89, BLN89, WL29);
sram_cell_6t_3 inst_cell_29_88 ( BL88, BLN88, WL29);
sram_cell_6t_3 inst_cell_29_87 ( BL87, BLN87, WL29);
sram_cell_6t_3 inst_cell_29_86 ( BL86, BLN86, WL29);
sram_cell_6t_3 inst_cell_29_85 ( BL85, BLN85, WL29);
sram_cell_6t_3 inst_cell_29_84 ( BL84, BLN84, WL29);
sram_cell_6t_3 inst_cell_29_83 ( BL83, BLN83, WL29);
sram_cell_6t_3 inst_cell_29_82 ( BL82, BLN82, WL29);
sram_cell_6t_3 inst_cell_29_81 ( BL81, BLN81, WL29);
sram_cell_6t_3 inst_cell_29_80 ( BL80, BLN80, WL29);
sram_cell_6t_3 inst_cell_29_79 ( BL79, BLN79, WL29);
sram_cell_6t_3 inst_cell_29_78 ( BL78, BLN78, WL29);
sram_cell_6t_3 inst_cell_29_77 ( BL77, BLN77, WL29);
sram_cell_6t_3 inst_cell_29_76 ( BL76, BLN76, WL29);
sram_cell_6t_3 inst_cell_29_75 ( BL75, BLN75, WL29);
sram_cell_6t_3 inst_cell_29_74 ( BL74, BLN74, WL29);
sram_cell_6t_3 inst_cell_29_73 ( BL73, BLN73, WL29);
sram_cell_6t_3 inst_cell_29_72 ( BL72, BLN72, WL29);
sram_cell_6t_3 inst_cell_29_71 ( BL71, BLN71, WL29);
sram_cell_6t_3 inst_cell_29_70 ( BL70, BLN70, WL29);
sram_cell_6t_3 inst_cell_29_69 ( BL69, BLN69, WL29);
sram_cell_6t_3 inst_cell_29_68 ( BL68, BLN68, WL29);
sram_cell_6t_3 inst_cell_29_67 ( BL67, BLN67, WL29);
sram_cell_6t_3 inst_cell_29_66 ( BL66, BLN66, WL29);
sram_cell_6t_3 inst_cell_29_65 ( BL65, BLN65, WL29);
sram_cell_6t_3 inst_cell_29_64 ( BL64, BLN64, WL29);
sram_cell_6t_3 inst_cell_29_63 ( BL63, BLN63, WL29);
sram_cell_6t_3 inst_cell_29_62 ( BL62, BLN62, WL29);
sram_cell_6t_3 inst_cell_29_61 ( BL61, BLN61, WL29);
sram_cell_6t_3 inst_cell_29_60 ( BL60, BLN60, WL29);
sram_cell_6t_3 inst_cell_29_59 ( BL59, BLN59, WL29);
sram_cell_6t_3 inst_cell_29_58 ( BL58, BLN58, WL29);
sram_cell_6t_3 inst_cell_29_57 ( BL57, BLN57, WL29);
sram_cell_6t_3 inst_cell_29_56 ( BL56, BLN56, WL29);
sram_cell_6t_3 inst_cell_29_55 ( BL55, BLN55, WL29);
sram_cell_6t_3 inst_cell_29_54 ( BL54, BLN54, WL29);
sram_cell_6t_3 inst_cell_29_53 ( BL53, BLN53, WL29);
sram_cell_6t_3 inst_cell_29_52 ( BL52, BLN52, WL29);
sram_cell_6t_3 inst_cell_29_51 ( BL51, BLN51, WL29);
sram_cell_6t_3 inst_cell_29_50 ( BL50, BLN50, WL29);
sram_cell_6t_3 inst_cell_29_49 ( BL49, BLN49, WL29);
sram_cell_6t_3 inst_cell_29_48 ( BL48, BLN48, WL29);
sram_cell_6t_3 inst_cell_29_47 ( BL47, BLN47, WL29);
sram_cell_6t_3 inst_cell_29_46 ( BL46, BLN46, WL29);
sram_cell_6t_3 inst_cell_29_45 ( BL45, BLN45, WL29);
sram_cell_6t_3 inst_cell_29_44 ( BL44, BLN44, WL29);
sram_cell_6t_3 inst_cell_29_43 ( BL43, BLN43, WL29);
sram_cell_6t_3 inst_cell_29_42 ( BL42, BLN42, WL29);
sram_cell_6t_3 inst_cell_29_41 ( BL41, BLN41, WL29);
sram_cell_6t_3 inst_cell_29_40 ( BL40, BLN40, WL29);
sram_cell_6t_3 inst_cell_29_39 ( BL39, BLN39, WL29);
sram_cell_6t_3 inst_cell_29_38 ( BL38, BLN38, WL29);
sram_cell_6t_3 inst_cell_29_37 ( BL37, BLN37, WL29);
sram_cell_6t_3 inst_cell_29_36 ( BL36, BLN36, WL29);
sram_cell_6t_3 inst_cell_29_35 ( BL35, BLN35, WL29);
sram_cell_6t_3 inst_cell_29_34 ( BL34, BLN34, WL29);
sram_cell_6t_3 inst_cell_29_33 ( BL33, BLN33, WL29);
sram_cell_6t_3 inst_cell_29_32 ( BL32, BLN32, WL29);
sram_cell_6t_3 inst_cell_29_31 ( BL31, BLN31, WL29);
sram_cell_6t_3 inst_cell_29_30 ( BL30, BLN30, WL29);
sram_cell_6t_3 inst_cell_29_29 ( BL29, BLN29, WL29);
sram_cell_6t_3 inst_cell_29_28 ( BL28, BLN28, WL29);
sram_cell_6t_3 inst_cell_29_27 ( BL27, BLN27, WL29);
sram_cell_6t_3 inst_cell_29_26 ( BL26, BLN26, WL29);
sram_cell_6t_3 inst_cell_29_25 ( BL25, BLN25, WL29);
sram_cell_6t_3 inst_cell_29_24 ( BL24, BLN24, WL29);
sram_cell_6t_3 inst_cell_29_23 ( BL23, BLN23, WL29);
sram_cell_6t_3 inst_cell_29_22 ( BL22, BLN22, WL29);
sram_cell_6t_3 inst_cell_29_21 ( BL21, BLN21, WL29);
sram_cell_6t_3 inst_cell_29_20 ( BL20, BLN20, WL29);
sram_cell_6t_3 inst_cell_29_19 ( BL19, BLN19, WL29);
sram_cell_6t_3 inst_cell_29_18 ( BL18, BLN18, WL29);
sram_cell_6t_3 inst_cell_29_17 ( BL17, BLN17, WL29);
sram_cell_6t_3 inst_cell_29_16 ( BL16, BLN16, WL29);
sram_cell_6t_3 inst_cell_29_15 ( BL15, BLN15, WL29);
sram_cell_6t_3 inst_cell_29_14 ( BL14, BLN14, WL29);
sram_cell_6t_3 inst_cell_29_13 ( BL13, BLN13, WL29);
sram_cell_6t_3 inst_cell_29_12 ( BL12, BLN12, WL29);
sram_cell_6t_3 inst_cell_29_11 ( BL11, BLN11, WL29);
sram_cell_6t_3 inst_cell_29_10 ( BL10, BLN10, WL29);
sram_cell_6t_3 inst_cell_29_9 ( BL9, BLN9, WL29);
sram_cell_6t_3 inst_cell_29_8 ( BL8, BLN8, WL29);
sram_cell_6t_3 inst_cell_29_7 ( BL7, BLN7, WL29);
sram_cell_6t_3 inst_cell_29_6 ( BL6, BLN6, WL29);
sram_cell_6t_3 inst_cell_29_5 ( BL5, BLN5, WL29);
sram_cell_6t_3 inst_cell_29_4 ( BL4, BLN4, WL29);
sram_cell_6t_3 inst_cell_29_3 ( BL3, BLN3, WL29);
sram_cell_6t_3 inst_cell_29_2 ( BL2, BLN2, WL29);
sram_cell_6t_3 inst_cell_29_1 ( BL1, BLN1, WL29);
sram_cell_6t_3 inst_cell_29_0 ( BL0, BLN0, WL29);
sram_cell_6t_3 inst_cell_28_127 ( BL127, BLN127, WL28);
sram_cell_6t_3 inst_cell_28_126 ( BL126, BLN126, WL28);
sram_cell_6t_3 inst_cell_28_125 ( BL125, BLN125, WL28);
sram_cell_6t_3 inst_cell_28_124 ( BL124, BLN124, WL28);
sram_cell_6t_3 inst_cell_28_123 ( BL123, BLN123, WL28);
sram_cell_6t_3 inst_cell_28_122 ( BL122, BLN122, WL28);
sram_cell_6t_3 inst_cell_28_121 ( BL121, BLN121, WL28);
sram_cell_6t_3 inst_cell_28_120 ( BL120, BLN120, WL28);
sram_cell_6t_3 inst_cell_28_119 ( BL119, BLN119, WL28);
sram_cell_6t_3 inst_cell_28_118 ( BL118, BLN118, WL28);
sram_cell_6t_3 inst_cell_28_117 ( BL117, BLN117, WL28);
sram_cell_6t_3 inst_cell_28_116 ( BL116, BLN116, WL28);
sram_cell_6t_3 inst_cell_28_115 ( BL115, BLN115, WL28);
sram_cell_6t_3 inst_cell_28_114 ( BL114, BLN114, WL28);
sram_cell_6t_3 inst_cell_28_113 ( BL113, BLN113, WL28);
sram_cell_6t_3 inst_cell_28_112 ( BL112, BLN112, WL28);
sram_cell_6t_3 inst_cell_28_111 ( BL111, BLN111, WL28);
sram_cell_6t_3 inst_cell_28_110 ( BL110, BLN110, WL28);
sram_cell_6t_3 inst_cell_28_109 ( BL109, BLN109, WL28);
sram_cell_6t_3 inst_cell_28_108 ( BL108, BLN108, WL28);
sram_cell_6t_3 inst_cell_28_107 ( BL107, BLN107, WL28);
sram_cell_6t_3 inst_cell_28_106 ( BL106, BLN106, WL28);
sram_cell_6t_3 inst_cell_28_105 ( BL105, BLN105, WL28);
sram_cell_6t_3 inst_cell_28_104 ( BL104, BLN104, WL28);
sram_cell_6t_3 inst_cell_28_103 ( BL103, BLN103, WL28);
sram_cell_6t_3 inst_cell_28_102 ( BL102, BLN102, WL28);
sram_cell_6t_3 inst_cell_28_101 ( BL101, BLN101, WL28);
sram_cell_6t_3 inst_cell_28_100 ( BL100, BLN100, WL28);
sram_cell_6t_3 inst_cell_28_99 ( BL99, BLN99, WL28);
sram_cell_6t_3 inst_cell_28_98 ( BL98, BLN98, WL28);
sram_cell_6t_3 inst_cell_28_97 ( BL97, BLN97, WL28);
sram_cell_6t_3 inst_cell_28_96 ( BL96, BLN96, WL28);
sram_cell_6t_3 inst_cell_28_95 ( BL95, BLN95, WL28);
sram_cell_6t_3 inst_cell_28_94 ( BL94, BLN94, WL28);
sram_cell_6t_3 inst_cell_28_93 ( BL93, BLN93, WL28);
sram_cell_6t_3 inst_cell_28_92 ( BL92, BLN92, WL28);
sram_cell_6t_3 inst_cell_28_91 ( BL91, BLN91, WL28);
sram_cell_6t_3 inst_cell_28_90 ( BL90, BLN90, WL28);
sram_cell_6t_3 inst_cell_28_89 ( BL89, BLN89, WL28);
sram_cell_6t_3 inst_cell_28_88 ( BL88, BLN88, WL28);
sram_cell_6t_3 inst_cell_28_87 ( BL87, BLN87, WL28);
sram_cell_6t_3 inst_cell_28_86 ( BL86, BLN86, WL28);
sram_cell_6t_3 inst_cell_28_85 ( BL85, BLN85, WL28);
sram_cell_6t_3 inst_cell_28_84 ( BL84, BLN84, WL28);
sram_cell_6t_3 inst_cell_28_83 ( BL83, BLN83, WL28);
sram_cell_6t_3 inst_cell_28_82 ( BL82, BLN82, WL28);
sram_cell_6t_3 inst_cell_28_81 ( BL81, BLN81, WL28);
sram_cell_6t_3 inst_cell_28_80 ( BL80, BLN80, WL28);
sram_cell_6t_3 inst_cell_28_79 ( BL79, BLN79, WL28);
sram_cell_6t_3 inst_cell_28_78 ( BL78, BLN78, WL28);
sram_cell_6t_3 inst_cell_28_77 ( BL77, BLN77, WL28);
sram_cell_6t_3 inst_cell_28_76 ( BL76, BLN76, WL28);
sram_cell_6t_3 inst_cell_28_75 ( BL75, BLN75, WL28);
sram_cell_6t_3 inst_cell_28_74 ( BL74, BLN74, WL28);
sram_cell_6t_3 inst_cell_28_73 ( BL73, BLN73, WL28);
sram_cell_6t_3 inst_cell_28_72 ( BL72, BLN72, WL28);
sram_cell_6t_3 inst_cell_28_71 ( BL71, BLN71, WL28);
sram_cell_6t_3 inst_cell_28_70 ( BL70, BLN70, WL28);
sram_cell_6t_3 inst_cell_28_69 ( BL69, BLN69, WL28);
sram_cell_6t_3 inst_cell_28_68 ( BL68, BLN68, WL28);
sram_cell_6t_3 inst_cell_28_67 ( BL67, BLN67, WL28);
sram_cell_6t_3 inst_cell_28_66 ( BL66, BLN66, WL28);
sram_cell_6t_3 inst_cell_28_65 ( BL65, BLN65, WL28);
sram_cell_6t_3 inst_cell_28_64 ( BL64, BLN64, WL28);
sram_cell_6t_3 inst_cell_28_63 ( BL63, BLN63, WL28);
sram_cell_6t_3 inst_cell_28_62 ( BL62, BLN62, WL28);
sram_cell_6t_3 inst_cell_28_61 ( BL61, BLN61, WL28);
sram_cell_6t_3 inst_cell_28_60 ( BL60, BLN60, WL28);
sram_cell_6t_3 inst_cell_28_59 ( BL59, BLN59, WL28);
sram_cell_6t_3 inst_cell_28_58 ( BL58, BLN58, WL28);
sram_cell_6t_3 inst_cell_28_57 ( BL57, BLN57, WL28);
sram_cell_6t_3 inst_cell_28_56 ( BL56, BLN56, WL28);
sram_cell_6t_3 inst_cell_28_55 ( BL55, BLN55, WL28);
sram_cell_6t_3 inst_cell_28_54 ( BL54, BLN54, WL28);
sram_cell_6t_3 inst_cell_28_53 ( BL53, BLN53, WL28);
sram_cell_6t_3 inst_cell_28_52 ( BL52, BLN52, WL28);
sram_cell_6t_3 inst_cell_28_51 ( BL51, BLN51, WL28);
sram_cell_6t_3 inst_cell_28_50 ( BL50, BLN50, WL28);
sram_cell_6t_3 inst_cell_28_49 ( BL49, BLN49, WL28);
sram_cell_6t_3 inst_cell_28_48 ( BL48, BLN48, WL28);
sram_cell_6t_3 inst_cell_28_47 ( BL47, BLN47, WL28);
sram_cell_6t_3 inst_cell_28_46 ( BL46, BLN46, WL28);
sram_cell_6t_3 inst_cell_28_45 ( BL45, BLN45, WL28);
sram_cell_6t_3 inst_cell_28_44 ( BL44, BLN44, WL28);
sram_cell_6t_3 inst_cell_28_43 ( BL43, BLN43, WL28);
sram_cell_6t_3 inst_cell_28_42 ( BL42, BLN42, WL28);
sram_cell_6t_3 inst_cell_28_41 ( BL41, BLN41, WL28);
sram_cell_6t_3 inst_cell_28_40 ( BL40, BLN40, WL28);
sram_cell_6t_3 inst_cell_28_39 ( BL39, BLN39, WL28);
sram_cell_6t_3 inst_cell_28_38 ( BL38, BLN38, WL28);
sram_cell_6t_3 inst_cell_28_37 ( BL37, BLN37, WL28);
sram_cell_6t_3 inst_cell_28_36 ( BL36, BLN36, WL28);
sram_cell_6t_3 inst_cell_28_35 ( BL35, BLN35, WL28);
sram_cell_6t_3 inst_cell_28_34 ( BL34, BLN34, WL28);
sram_cell_6t_3 inst_cell_28_33 ( BL33, BLN33, WL28);
sram_cell_6t_3 inst_cell_28_32 ( BL32, BLN32, WL28);
sram_cell_6t_3 inst_cell_28_31 ( BL31, BLN31, WL28);
sram_cell_6t_3 inst_cell_28_30 ( BL30, BLN30, WL28);
sram_cell_6t_3 inst_cell_28_29 ( BL29, BLN29, WL28);
sram_cell_6t_3 inst_cell_28_28 ( BL28, BLN28, WL28);
sram_cell_6t_3 inst_cell_28_27 ( BL27, BLN27, WL28);
sram_cell_6t_3 inst_cell_28_26 ( BL26, BLN26, WL28);
sram_cell_6t_3 inst_cell_28_25 ( BL25, BLN25, WL28);
sram_cell_6t_3 inst_cell_28_24 ( BL24, BLN24, WL28);
sram_cell_6t_3 inst_cell_28_23 ( BL23, BLN23, WL28);
sram_cell_6t_3 inst_cell_28_22 ( BL22, BLN22, WL28);
sram_cell_6t_3 inst_cell_28_21 ( BL21, BLN21, WL28);
sram_cell_6t_3 inst_cell_28_20 ( BL20, BLN20, WL28);
sram_cell_6t_3 inst_cell_28_19 ( BL19, BLN19, WL28);
sram_cell_6t_3 inst_cell_28_18 ( BL18, BLN18, WL28);
sram_cell_6t_3 inst_cell_28_17 ( BL17, BLN17, WL28);
sram_cell_6t_3 inst_cell_28_16 ( BL16, BLN16, WL28);
sram_cell_6t_3 inst_cell_28_15 ( BL15, BLN15, WL28);
sram_cell_6t_3 inst_cell_28_14 ( BL14, BLN14, WL28);
sram_cell_6t_3 inst_cell_28_13 ( BL13, BLN13, WL28);
sram_cell_6t_3 inst_cell_28_12 ( BL12, BLN12, WL28);
sram_cell_6t_3 inst_cell_28_11 ( BL11, BLN11, WL28);
sram_cell_6t_3 inst_cell_28_10 ( BL10, BLN10, WL28);
sram_cell_6t_3 inst_cell_28_9 ( BL9, BLN9, WL28);
sram_cell_6t_3 inst_cell_28_8 ( BL8, BLN8, WL28);
sram_cell_6t_3 inst_cell_28_7 ( BL7, BLN7, WL28);
sram_cell_6t_3 inst_cell_28_6 ( BL6, BLN6, WL28);
sram_cell_6t_3 inst_cell_28_5 ( BL5, BLN5, WL28);
sram_cell_6t_3 inst_cell_28_4 ( BL4, BLN4, WL28);
sram_cell_6t_3 inst_cell_28_3 ( BL3, BLN3, WL28);
sram_cell_6t_3 inst_cell_28_2 ( BL2, BLN2, WL28);
sram_cell_6t_3 inst_cell_28_1 ( BL1, BLN1, WL28);
sram_cell_6t_3 inst_cell_28_0 ( BL0, BLN0, WL28);
sram_cell_6t_3 inst_cell_27_127 ( BL127, BLN127, WL27);
sram_cell_6t_3 inst_cell_27_126 ( BL126, BLN126, WL27);
sram_cell_6t_3 inst_cell_27_125 ( BL125, BLN125, WL27);
sram_cell_6t_3 inst_cell_27_124 ( BL124, BLN124, WL27);
sram_cell_6t_3 inst_cell_27_123 ( BL123, BLN123, WL27);
sram_cell_6t_3 inst_cell_27_122 ( BL122, BLN122, WL27);
sram_cell_6t_3 inst_cell_27_121 ( BL121, BLN121, WL27);
sram_cell_6t_3 inst_cell_27_120 ( BL120, BLN120, WL27);
sram_cell_6t_3 inst_cell_27_119 ( BL119, BLN119, WL27);
sram_cell_6t_3 inst_cell_27_118 ( BL118, BLN118, WL27);
sram_cell_6t_3 inst_cell_27_117 ( BL117, BLN117, WL27);
sram_cell_6t_3 inst_cell_27_116 ( BL116, BLN116, WL27);
sram_cell_6t_3 inst_cell_27_115 ( BL115, BLN115, WL27);
sram_cell_6t_3 inst_cell_27_114 ( BL114, BLN114, WL27);
sram_cell_6t_3 inst_cell_27_113 ( BL113, BLN113, WL27);
sram_cell_6t_3 inst_cell_27_112 ( BL112, BLN112, WL27);
sram_cell_6t_3 inst_cell_27_111 ( BL111, BLN111, WL27);
sram_cell_6t_3 inst_cell_27_110 ( BL110, BLN110, WL27);
sram_cell_6t_3 inst_cell_27_109 ( BL109, BLN109, WL27);
sram_cell_6t_3 inst_cell_27_108 ( BL108, BLN108, WL27);
sram_cell_6t_3 inst_cell_27_107 ( BL107, BLN107, WL27);
sram_cell_6t_3 inst_cell_27_106 ( BL106, BLN106, WL27);
sram_cell_6t_3 inst_cell_27_105 ( BL105, BLN105, WL27);
sram_cell_6t_3 inst_cell_27_104 ( BL104, BLN104, WL27);
sram_cell_6t_3 inst_cell_27_103 ( BL103, BLN103, WL27);
sram_cell_6t_3 inst_cell_27_102 ( BL102, BLN102, WL27);
sram_cell_6t_3 inst_cell_27_101 ( BL101, BLN101, WL27);
sram_cell_6t_3 inst_cell_27_100 ( BL100, BLN100, WL27);
sram_cell_6t_3 inst_cell_27_99 ( BL99, BLN99, WL27);
sram_cell_6t_3 inst_cell_27_98 ( BL98, BLN98, WL27);
sram_cell_6t_3 inst_cell_27_97 ( BL97, BLN97, WL27);
sram_cell_6t_3 inst_cell_27_96 ( BL96, BLN96, WL27);
sram_cell_6t_3 inst_cell_27_95 ( BL95, BLN95, WL27);
sram_cell_6t_3 inst_cell_27_94 ( BL94, BLN94, WL27);
sram_cell_6t_3 inst_cell_27_93 ( BL93, BLN93, WL27);
sram_cell_6t_3 inst_cell_27_92 ( BL92, BLN92, WL27);
sram_cell_6t_3 inst_cell_27_91 ( BL91, BLN91, WL27);
sram_cell_6t_3 inst_cell_27_90 ( BL90, BLN90, WL27);
sram_cell_6t_3 inst_cell_27_89 ( BL89, BLN89, WL27);
sram_cell_6t_3 inst_cell_27_88 ( BL88, BLN88, WL27);
sram_cell_6t_3 inst_cell_27_87 ( BL87, BLN87, WL27);
sram_cell_6t_3 inst_cell_27_86 ( BL86, BLN86, WL27);
sram_cell_6t_3 inst_cell_27_85 ( BL85, BLN85, WL27);
sram_cell_6t_3 inst_cell_27_84 ( BL84, BLN84, WL27);
sram_cell_6t_3 inst_cell_27_83 ( BL83, BLN83, WL27);
sram_cell_6t_3 inst_cell_27_82 ( BL82, BLN82, WL27);
sram_cell_6t_3 inst_cell_27_81 ( BL81, BLN81, WL27);
sram_cell_6t_3 inst_cell_27_80 ( BL80, BLN80, WL27);
sram_cell_6t_3 inst_cell_27_79 ( BL79, BLN79, WL27);
sram_cell_6t_3 inst_cell_27_78 ( BL78, BLN78, WL27);
sram_cell_6t_3 inst_cell_27_77 ( BL77, BLN77, WL27);
sram_cell_6t_3 inst_cell_27_76 ( BL76, BLN76, WL27);
sram_cell_6t_3 inst_cell_27_75 ( BL75, BLN75, WL27);
sram_cell_6t_3 inst_cell_27_74 ( BL74, BLN74, WL27);
sram_cell_6t_3 inst_cell_27_73 ( BL73, BLN73, WL27);
sram_cell_6t_3 inst_cell_27_72 ( BL72, BLN72, WL27);
sram_cell_6t_3 inst_cell_27_71 ( BL71, BLN71, WL27);
sram_cell_6t_3 inst_cell_27_70 ( BL70, BLN70, WL27);
sram_cell_6t_3 inst_cell_27_69 ( BL69, BLN69, WL27);
sram_cell_6t_3 inst_cell_27_68 ( BL68, BLN68, WL27);
sram_cell_6t_3 inst_cell_27_67 ( BL67, BLN67, WL27);
sram_cell_6t_3 inst_cell_27_66 ( BL66, BLN66, WL27);
sram_cell_6t_3 inst_cell_27_65 ( BL65, BLN65, WL27);
sram_cell_6t_3 inst_cell_27_64 ( BL64, BLN64, WL27);
sram_cell_6t_3 inst_cell_27_63 ( BL63, BLN63, WL27);
sram_cell_6t_3 inst_cell_27_62 ( BL62, BLN62, WL27);
sram_cell_6t_3 inst_cell_27_61 ( BL61, BLN61, WL27);
sram_cell_6t_3 inst_cell_27_60 ( BL60, BLN60, WL27);
sram_cell_6t_3 inst_cell_27_59 ( BL59, BLN59, WL27);
sram_cell_6t_3 inst_cell_27_58 ( BL58, BLN58, WL27);
sram_cell_6t_3 inst_cell_27_57 ( BL57, BLN57, WL27);
sram_cell_6t_3 inst_cell_27_56 ( BL56, BLN56, WL27);
sram_cell_6t_3 inst_cell_27_55 ( BL55, BLN55, WL27);
sram_cell_6t_3 inst_cell_27_54 ( BL54, BLN54, WL27);
sram_cell_6t_3 inst_cell_27_53 ( BL53, BLN53, WL27);
sram_cell_6t_3 inst_cell_27_52 ( BL52, BLN52, WL27);
sram_cell_6t_3 inst_cell_27_51 ( BL51, BLN51, WL27);
sram_cell_6t_3 inst_cell_27_50 ( BL50, BLN50, WL27);
sram_cell_6t_3 inst_cell_27_49 ( BL49, BLN49, WL27);
sram_cell_6t_3 inst_cell_27_48 ( BL48, BLN48, WL27);
sram_cell_6t_3 inst_cell_27_47 ( BL47, BLN47, WL27);
sram_cell_6t_3 inst_cell_27_46 ( BL46, BLN46, WL27);
sram_cell_6t_3 inst_cell_27_45 ( BL45, BLN45, WL27);
sram_cell_6t_3 inst_cell_27_44 ( BL44, BLN44, WL27);
sram_cell_6t_3 inst_cell_27_43 ( BL43, BLN43, WL27);
sram_cell_6t_3 inst_cell_27_42 ( BL42, BLN42, WL27);
sram_cell_6t_3 inst_cell_27_41 ( BL41, BLN41, WL27);
sram_cell_6t_3 inst_cell_27_40 ( BL40, BLN40, WL27);
sram_cell_6t_3 inst_cell_27_39 ( BL39, BLN39, WL27);
sram_cell_6t_3 inst_cell_27_38 ( BL38, BLN38, WL27);
sram_cell_6t_3 inst_cell_27_37 ( BL37, BLN37, WL27);
sram_cell_6t_3 inst_cell_27_36 ( BL36, BLN36, WL27);
sram_cell_6t_3 inst_cell_27_35 ( BL35, BLN35, WL27);
sram_cell_6t_3 inst_cell_27_34 ( BL34, BLN34, WL27);
sram_cell_6t_3 inst_cell_27_33 ( BL33, BLN33, WL27);
sram_cell_6t_3 inst_cell_27_32 ( BL32, BLN32, WL27);
sram_cell_6t_3 inst_cell_27_31 ( BL31, BLN31, WL27);
sram_cell_6t_3 inst_cell_27_30 ( BL30, BLN30, WL27);
sram_cell_6t_3 inst_cell_27_29 ( BL29, BLN29, WL27);
sram_cell_6t_3 inst_cell_27_28 ( BL28, BLN28, WL27);
sram_cell_6t_3 inst_cell_27_27 ( BL27, BLN27, WL27);
sram_cell_6t_3 inst_cell_27_26 ( BL26, BLN26, WL27);
sram_cell_6t_3 inst_cell_27_25 ( BL25, BLN25, WL27);
sram_cell_6t_3 inst_cell_27_24 ( BL24, BLN24, WL27);
sram_cell_6t_3 inst_cell_27_23 ( BL23, BLN23, WL27);
sram_cell_6t_3 inst_cell_27_22 ( BL22, BLN22, WL27);
sram_cell_6t_3 inst_cell_27_21 ( BL21, BLN21, WL27);
sram_cell_6t_3 inst_cell_27_20 ( BL20, BLN20, WL27);
sram_cell_6t_3 inst_cell_27_19 ( BL19, BLN19, WL27);
sram_cell_6t_3 inst_cell_27_18 ( BL18, BLN18, WL27);
sram_cell_6t_3 inst_cell_27_17 ( BL17, BLN17, WL27);
sram_cell_6t_3 inst_cell_27_16 ( BL16, BLN16, WL27);
sram_cell_6t_3 inst_cell_27_15 ( BL15, BLN15, WL27);
sram_cell_6t_3 inst_cell_27_14 ( BL14, BLN14, WL27);
sram_cell_6t_3 inst_cell_27_13 ( BL13, BLN13, WL27);
sram_cell_6t_3 inst_cell_27_12 ( BL12, BLN12, WL27);
sram_cell_6t_3 inst_cell_27_11 ( BL11, BLN11, WL27);
sram_cell_6t_3 inst_cell_27_10 ( BL10, BLN10, WL27);
sram_cell_6t_3 inst_cell_27_9 ( BL9, BLN9, WL27);
sram_cell_6t_3 inst_cell_27_8 ( BL8, BLN8, WL27);
sram_cell_6t_3 inst_cell_27_7 ( BL7, BLN7, WL27);
sram_cell_6t_3 inst_cell_27_6 ( BL6, BLN6, WL27);
sram_cell_6t_3 inst_cell_27_5 ( BL5, BLN5, WL27);
sram_cell_6t_3 inst_cell_27_4 ( BL4, BLN4, WL27);
sram_cell_6t_3 inst_cell_27_3 ( BL3, BLN3, WL27);
sram_cell_6t_3 inst_cell_27_2 ( BL2, BLN2, WL27);
sram_cell_6t_3 inst_cell_27_1 ( BL1, BLN1, WL27);
sram_cell_6t_3 inst_cell_27_0 ( BL0, BLN0, WL27);
sram_cell_6t_3 inst_cell_26_127 ( BL127, BLN127, WL26);
sram_cell_6t_3 inst_cell_26_126 ( BL126, BLN126, WL26);
sram_cell_6t_3 inst_cell_26_125 ( BL125, BLN125, WL26);
sram_cell_6t_3 inst_cell_26_124 ( BL124, BLN124, WL26);
sram_cell_6t_3 inst_cell_26_123 ( BL123, BLN123, WL26);
sram_cell_6t_3 inst_cell_26_122 ( BL122, BLN122, WL26);
sram_cell_6t_3 inst_cell_26_121 ( BL121, BLN121, WL26);
sram_cell_6t_3 inst_cell_26_120 ( BL120, BLN120, WL26);
sram_cell_6t_3 inst_cell_26_119 ( BL119, BLN119, WL26);
sram_cell_6t_3 inst_cell_26_118 ( BL118, BLN118, WL26);
sram_cell_6t_3 inst_cell_26_117 ( BL117, BLN117, WL26);
sram_cell_6t_3 inst_cell_26_116 ( BL116, BLN116, WL26);
sram_cell_6t_3 inst_cell_26_115 ( BL115, BLN115, WL26);
sram_cell_6t_3 inst_cell_26_114 ( BL114, BLN114, WL26);
sram_cell_6t_3 inst_cell_26_113 ( BL113, BLN113, WL26);
sram_cell_6t_3 inst_cell_26_112 ( BL112, BLN112, WL26);
sram_cell_6t_3 inst_cell_26_111 ( BL111, BLN111, WL26);
sram_cell_6t_3 inst_cell_26_110 ( BL110, BLN110, WL26);
sram_cell_6t_3 inst_cell_26_109 ( BL109, BLN109, WL26);
sram_cell_6t_3 inst_cell_26_108 ( BL108, BLN108, WL26);
sram_cell_6t_3 inst_cell_26_107 ( BL107, BLN107, WL26);
sram_cell_6t_3 inst_cell_26_106 ( BL106, BLN106, WL26);
sram_cell_6t_3 inst_cell_26_105 ( BL105, BLN105, WL26);
sram_cell_6t_3 inst_cell_26_104 ( BL104, BLN104, WL26);
sram_cell_6t_3 inst_cell_26_103 ( BL103, BLN103, WL26);
sram_cell_6t_3 inst_cell_26_102 ( BL102, BLN102, WL26);
sram_cell_6t_3 inst_cell_26_101 ( BL101, BLN101, WL26);
sram_cell_6t_3 inst_cell_26_100 ( BL100, BLN100, WL26);
sram_cell_6t_3 inst_cell_26_99 ( BL99, BLN99, WL26);
sram_cell_6t_3 inst_cell_26_98 ( BL98, BLN98, WL26);
sram_cell_6t_3 inst_cell_26_97 ( BL97, BLN97, WL26);
sram_cell_6t_3 inst_cell_26_96 ( BL96, BLN96, WL26);
sram_cell_6t_3 inst_cell_26_95 ( BL95, BLN95, WL26);
sram_cell_6t_3 inst_cell_26_94 ( BL94, BLN94, WL26);
sram_cell_6t_3 inst_cell_26_93 ( BL93, BLN93, WL26);
sram_cell_6t_3 inst_cell_26_92 ( BL92, BLN92, WL26);
sram_cell_6t_3 inst_cell_26_91 ( BL91, BLN91, WL26);
sram_cell_6t_3 inst_cell_26_90 ( BL90, BLN90, WL26);
sram_cell_6t_3 inst_cell_26_89 ( BL89, BLN89, WL26);
sram_cell_6t_3 inst_cell_26_88 ( BL88, BLN88, WL26);
sram_cell_6t_3 inst_cell_26_87 ( BL87, BLN87, WL26);
sram_cell_6t_3 inst_cell_26_86 ( BL86, BLN86, WL26);
sram_cell_6t_3 inst_cell_26_85 ( BL85, BLN85, WL26);
sram_cell_6t_3 inst_cell_26_84 ( BL84, BLN84, WL26);
sram_cell_6t_3 inst_cell_26_83 ( BL83, BLN83, WL26);
sram_cell_6t_3 inst_cell_26_82 ( BL82, BLN82, WL26);
sram_cell_6t_3 inst_cell_26_81 ( BL81, BLN81, WL26);
sram_cell_6t_3 inst_cell_26_80 ( BL80, BLN80, WL26);
sram_cell_6t_3 inst_cell_26_79 ( BL79, BLN79, WL26);
sram_cell_6t_3 inst_cell_26_78 ( BL78, BLN78, WL26);
sram_cell_6t_3 inst_cell_26_77 ( BL77, BLN77, WL26);
sram_cell_6t_3 inst_cell_26_76 ( BL76, BLN76, WL26);
sram_cell_6t_3 inst_cell_26_75 ( BL75, BLN75, WL26);
sram_cell_6t_3 inst_cell_26_74 ( BL74, BLN74, WL26);
sram_cell_6t_3 inst_cell_26_73 ( BL73, BLN73, WL26);
sram_cell_6t_3 inst_cell_26_72 ( BL72, BLN72, WL26);
sram_cell_6t_3 inst_cell_26_71 ( BL71, BLN71, WL26);
sram_cell_6t_3 inst_cell_26_70 ( BL70, BLN70, WL26);
sram_cell_6t_3 inst_cell_26_69 ( BL69, BLN69, WL26);
sram_cell_6t_3 inst_cell_26_68 ( BL68, BLN68, WL26);
sram_cell_6t_3 inst_cell_26_67 ( BL67, BLN67, WL26);
sram_cell_6t_3 inst_cell_26_66 ( BL66, BLN66, WL26);
sram_cell_6t_3 inst_cell_26_65 ( BL65, BLN65, WL26);
sram_cell_6t_3 inst_cell_26_64 ( BL64, BLN64, WL26);
sram_cell_6t_3 inst_cell_26_63 ( BL63, BLN63, WL26);
sram_cell_6t_3 inst_cell_26_62 ( BL62, BLN62, WL26);
sram_cell_6t_3 inst_cell_26_61 ( BL61, BLN61, WL26);
sram_cell_6t_3 inst_cell_26_60 ( BL60, BLN60, WL26);
sram_cell_6t_3 inst_cell_26_59 ( BL59, BLN59, WL26);
sram_cell_6t_3 inst_cell_26_58 ( BL58, BLN58, WL26);
sram_cell_6t_3 inst_cell_26_57 ( BL57, BLN57, WL26);
sram_cell_6t_3 inst_cell_26_56 ( BL56, BLN56, WL26);
sram_cell_6t_3 inst_cell_26_55 ( BL55, BLN55, WL26);
sram_cell_6t_3 inst_cell_26_54 ( BL54, BLN54, WL26);
sram_cell_6t_3 inst_cell_26_53 ( BL53, BLN53, WL26);
sram_cell_6t_3 inst_cell_26_52 ( BL52, BLN52, WL26);
sram_cell_6t_3 inst_cell_26_51 ( BL51, BLN51, WL26);
sram_cell_6t_3 inst_cell_26_50 ( BL50, BLN50, WL26);
sram_cell_6t_3 inst_cell_26_49 ( BL49, BLN49, WL26);
sram_cell_6t_3 inst_cell_26_48 ( BL48, BLN48, WL26);
sram_cell_6t_3 inst_cell_26_47 ( BL47, BLN47, WL26);
sram_cell_6t_3 inst_cell_26_46 ( BL46, BLN46, WL26);
sram_cell_6t_3 inst_cell_26_45 ( BL45, BLN45, WL26);
sram_cell_6t_3 inst_cell_26_44 ( BL44, BLN44, WL26);
sram_cell_6t_3 inst_cell_26_43 ( BL43, BLN43, WL26);
sram_cell_6t_3 inst_cell_26_42 ( BL42, BLN42, WL26);
sram_cell_6t_3 inst_cell_26_41 ( BL41, BLN41, WL26);
sram_cell_6t_3 inst_cell_26_40 ( BL40, BLN40, WL26);
sram_cell_6t_3 inst_cell_26_39 ( BL39, BLN39, WL26);
sram_cell_6t_3 inst_cell_26_38 ( BL38, BLN38, WL26);
sram_cell_6t_3 inst_cell_26_37 ( BL37, BLN37, WL26);
sram_cell_6t_3 inst_cell_26_36 ( BL36, BLN36, WL26);
sram_cell_6t_3 inst_cell_26_35 ( BL35, BLN35, WL26);
sram_cell_6t_3 inst_cell_26_34 ( BL34, BLN34, WL26);
sram_cell_6t_3 inst_cell_26_33 ( BL33, BLN33, WL26);
sram_cell_6t_3 inst_cell_26_32 ( BL32, BLN32, WL26);
sram_cell_6t_3 inst_cell_26_31 ( BL31, BLN31, WL26);
sram_cell_6t_3 inst_cell_26_30 ( BL30, BLN30, WL26);
sram_cell_6t_3 inst_cell_26_29 ( BL29, BLN29, WL26);
sram_cell_6t_3 inst_cell_26_28 ( BL28, BLN28, WL26);
sram_cell_6t_3 inst_cell_26_27 ( BL27, BLN27, WL26);
sram_cell_6t_3 inst_cell_26_26 ( BL26, BLN26, WL26);
sram_cell_6t_3 inst_cell_26_25 ( BL25, BLN25, WL26);
sram_cell_6t_3 inst_cell_26_24 ( BL24, BLN24, WL26);
sram_cell_6t_3 inst_cell_26_23 ( BL23, BLN23, WL26);
sram_cell_6t_3 inst_cell_26_22 ( BL22, BLN22, WL26);
sram_cell_6t_3 inst_cell_26_21 ( BL21, BLN21, WL26);
sram_cell_6t_3 inst_cell_26_20 ( BL20, BLN20, WL26);
sram_cell_6t_3 inst_cell_26_19 ( BL19, BLN19, WL26);
sram_cell_6t_3 inst_cell_26_18 ( BL18, BLN18, WL26);
sram_cell_6t_3 inst_cell_26_17 ( BL17, BLN17, WL26);
sram_cell_6t_3 inst_cell_26_16 ( BL16, BLN16, WL26);
sram_cell_6t_3 inst_cell_26_15 ( BL15, BLN15, WL26);
sram_cell_6t_3 inst_cell_26_14 ( BL14, BLN14, WL26);
sram_cell_6t_3 inst_cell_26_13 ( BL13, BLN13, WL26);
sram_cell_6t_3 inst_cell_26_12 ( BL12, BLN12, WL26);
sram_cell_6t_3 inst_cell_26_11 ( BL11, BLN11, WL26);
sram_cell_6t_3 inst_cell_26_10 ( BL10, BLN10, WL26);
sram_cell_6t_3 inst_cell_26_9 ( BL9, BLN9, WL26);
sram_cell_6t_3 inst_cell_26_8 ( BL8, BLN8, WL26);
sram_cell_6t_3 inst_cell_26_7 ( BL7, BLN7, WL26);
sram_cell_6t_3 inst_cell_26_6 ( BL6, BLN6, WL26);
sram_cell_6t_3 inst_cell_26_5 ( BL5, BLN5, WL26);
sram_cell_6t_3 inst_cell_26_4 ( BL4, BLN4, WL26);
sram_cell_6t_3 inst_cell_26_3 ( BL3, BLN3, WL26);
sram_cell_6t_3 inst_cell_26_2 ( BL2, BLN2, WL26);
sram_cell_6t_3 inst_cell_26_1 ( BL1, BLN1, WL26);
sram_cell_6t_3 inst_cell_26_0 ( BL0, BLN0, WL26);
sram_cell_6t_3 inst_cell_25_127 ( BL127, BLN127, WL25);
sram_cell_6t_3 inst_cell_25_126 ( BL126, BLN126, WL25);
sram_cell_6t_3 inst_cell_25_125 ( BL125, BLN125, WL25);
sram_cell_6t_3 inst_cell_25_124 ( BL124, BLN124, WL25);
sram_cell_6t_3 inst_cell_25_123 ( BL123, BLN123, WL25);
sram_cell_6t_3 inst_cell_25_122 ( BL122, BLN122, WL25);
sram_cell_6t_3 inst_cell_25_121 ( BL121, BLN121, WL25);
sram_cell_6t_3 inst_cell_25_120 ( BL120, BLN120, WL25);
sram_cell_6t_3 inst_cell_25_119 ( BL119, BLN119, WL25);
sram_cell_6t_3 inst_cell_25_118 ( BL118, BLN118, WL25);
sram_cell_6t_3 inst_cell_25_117 ( BL117, BLN117, WL25);
sram_cell_6t_3 inst_cell_25_116 ( BL116, BLN116, WL25);
sram_cell_6t_3 inst_cell_25_115 ( BL115, BLN115, WL25);
sram_cell_6t_3 inst_cell_25_114 ( BL114, BLN114, WL25);
sram_cell_6t_3 inst_cell_25_113 ( BL113, BLN113, WL25);
sram_cell_6t_3 inst_cell_25_112 ( BL112, BLN112, WL25);
sram_cell_6t_3 inst_cell_25_111 ( BL111, BLN111, WL25);
sram_cell_6t_3 inst_cell_25_110 ( BL110, BLN110, WL25);
sram_cell_6t_3 inst_cell_25_109 ( BL109, BLN109, WL25);
sram_cell_6t_3 inst_cell_25_108 ( BL108, BLN108, WL25);
sram_cell_6t_3 inst_cell_25_107 ( BL107, BLN107, WL25);
sram_cell_6t_3 inst_cell_25_106 ( BL106, BLN106, WL25);
sram_cell_6t_3 inst_cell_25_105 ( BL105, BLN105, WL25);
sram_cell_6t_3 inst_cell_25_104 ( BL104, BLN104, WL25);
sram_cell_6t_3 inst_cell_25_103 ( BL103, BLN103, WL25);
sram_cell_6t_3 inst_cell_25_102 ( BL102, BLN102, WL25);
sram_cell_6t_3 inst_cell_25_101 ( BL101, BLN101, WL25);
sram_cell_6t_3 inst_cell_25_100 ( BL100, BLN100, WL25);
sram_cell_6t_3 inst_cell_25_99 ( BL99, BLN99, WL25);
sram_cell_6t_3 inst_cell_25_98 ( BL98, BLN98, WL25);
sram_cell_6t_3 inst_cell_25_97 ( BL97, BLN97, WL25);
sram_cell_6t_3 inst_cell_25_96 ( BL96, BLN96, WL25);
sram_cell_6t_3 inst_cell_25_95 ( BL95, BLN95, WL25);
sram_cell_6t_3 inst_cell_25_94 ( BL94, BLN94, WL25);
sram_cell_6t_3 inst_cell_25_93 ( BL93, BLN93, WL25);
sram_cell_6t_3 inst_cell_25_92 ( BL92, BLN92, WL25);
sram_cell_6t_3 inst_cell_25_91 ( BL91, BLN91, WL25);
sram_cell_6t_3 inst_cell_25_90 ( BL90, BLN90, WL25);
sram_cell_6t_3 inst_cell_25_89 ( BL89, BLN89, WL25);
sram_cell_6t_3 inst_cell_25_88 ( BL88, BLN88, WL25);
sram_cell_6t_3 inst_cell_25_87 ( BL87, BLN87, WL25);
sram_cell_6t_3 inst_cell_25_86 ( BL86, BLN86, WL25);
sram_cell_6t_3 inst_cell_25_85 ( BL85, BLN85, WL25);
sram_cell_6t_3 inst_cell_25_84 ( BL84, BLN84, WL25);
sram_cell_6t_3 inst_cell_25_83 ( BL83, BLN83, WL25);
sram_cell_6t_3 inst_cell_25_82 ( BL82, BLN82, WL25);
sram_cell_6t_3 inst_cell_25_81 ( BL81, BLN81, WL25);
sram_cell_6t_3 inst_cell_25_80 ( BL80, BLN80, WL25);
sram_cell_6t_3 inst_cell_25_79 ( BL79, BLN79, WL25);
sram_cell_6t_3 inst_cell_25_78 ( BL78, BLN78, WL25);
sram_cell_6t_3 inst_cell_25_77 ( BL77, BLN77, WL25);
sram_cell_6t_3 inst_cell_25_76 ( BL76, BLN76, WL25);
sram_cell_6t_3 inst_cell_25_75 ( BL75, BLN75, WL25);
sram_cell_6t_3 inst_cell_25_74 ( BL74, BLN74, WL25);
sram_cell_6t_3 inst_cell_25_73 ( BL73, BLN73, WL25);
sram_cell_6t_3 inst_cell_25_72 ( BL72, BLN72, WL25);
sram_cell_6t_3 inst_cell_25_71 ( BL71, BLN71, WL25);
sram_cell_6t_3 inst_cell_25_70 ( BL70, BLN70, WL25);
sram_cell_6t_3 inst_cell_25_69 ( BL69, BLN69, WL25);
sram_cell_6t_3 inst_cell_25_68 ( BL68, BLN68, WL25);
sram_cell_6t_3 inst_cell_25_67 ( BL67, BLN67, WL25);
sram_cell_6t_3 inst_cell_25_66 ( BL66, BLN66, WL25);
sram_cell_6t_3 inst_cell_25_65 ( BL65, BLN65, WL25);
sram_cell_6t_3 inst_cell_25_64 ( BL64, BLN64, WL25);
sram_cell_6t_3 inst_cell_25_63 ( BL63, BLN63, WL25);
sram_cell_6t_3 inst_cell_25_62 ( BL62, BLN62, WL25);
sram_cell_6t_3 inst_cell_25_61 ( BL61, BLN61, WL25);
sram_cell_6t_3 inst_cell_25_60 ( BL60, BLN60, WL25);
sram_cell_6t_3 inst_cell_25_59 ( BL59, BLN59, WL25);
sram_cell_6t_3 inst_cell_25_58 ( BL58, BLN58, WL25);
sram_cell_6t_3 inst_cell_25_57 ( BL57, BLN57, WL25);
sram_cell_6t_3 inst_cell_25_56 ( BL56, BLN56, WL25);
sram_cell_6t_3 inst_cell_25_55 ( BL55, BLN55, WL25);
sram_cell_6t_3 inst_cell_25_54 ( BL54, BLN54, WL25);
sram_cell_6t_3 inst_cell_25_53 ( BL53, BLN53, WL25);
sram_cell_6t_3 inst_cell_25_52 ( BL52, BLN52, WL25);
sram_cell_6t_3 inst_cell_25_51 ( BL51, BLN51, WL25);
sram_cell_6t_3 inst_cell_25_50 ( BL50, BLN50, WL25);
sram_cell_6t_3 inst_cell_25_49 ( BL49, BLN49, WL25);
sram_cell_6t_3 inst_cell_25_48 ( BL48, BLN48, WL25);
sram_cell_6t_3 inst_cell_25_47 ( BL47, BLN47, WL25);
sram_cell_6t_3 inst_cell_25_46 ( BL46, BLN46, WL25);
sram_cell_6t_3 inst_cell_25_45 ( BL45, BLN45, WL25);
sram_cell_6t_3 inst_cell_25_44 ( BL44, BLN44, WL25);
sram_cell_6t_3 inst_cell_25_43 ( BL43, BLN43, WL25);
sram_cell_6t_3 inst_cell_25_42 ( BL42, BLN42, WL25);
sram_cell_6t_3 inst_cell_25_41 ( BL41, BLN41, WL25);
sram_cell_6t_3 inst_cell_25_40 ( BL40, BLN40, WL25);
sram_cell_6t_3 inst_cell_25_39 ( BL39, BLN39, WL25);
sram_cell_6t_3 inst_cell_25_38 ( BL38, BLN38, WL25);
sram_cell_6t_3 inst_cell_25_37 ( BL37, BLN37, WL25);
sram_cell_6t_3 inst_cell_25_36 ( BL36, BLN36, WL25);
sram_cell_6t_3 inst_cell_25_35 ( BL35, BLN35, WL25);
sram_cell_6t_3 inst_cell_25_34 ( BL34, BLN34, WL25);
sram_cell_6t_3 inst_cell_25_33 ( BL33, BLN33, WL25);
sram_cell_6t_3 inst_cell_25_32 ( BL32, BLN32, WL25);
sram_cell_6t_3 inst_cell_25_31 ( BL31, BLN31, WL25);
sram_cell_6t_3 inst_cell_25_30 ( BL30, BLN30, WL25);
sram_cell_6t_3 inst_cell_25_29 ( BL29, BLN29, WL25);
sram_cell_6t_3 inst_cell_25_28 ( BL28, BLN28, WL25);
sram_cell_6t_3 inst_cell_25_27 ( BL27, BLN27, WL25);
sram_cell_6t_3 inst_cell_25_26 ( BL26, BLN26, WL25);
sram_cell_6t_3 inst_cell_25_25 ( BL25, BLN25, WL25);
sram_cell_6t_3 inst_cell_25_24 ( BL24, BLN24, WL25);
sram_cell_6t_3 inst_cell_25_23 ( BL23, BLN23, WL25);
sram_cell_6t_3 inst_cell_25_22 ( BL22, BLN22, WL25);
sram_cell_6t_3 inst_cell_25_21 ( BL21, BLN21, WL25);
sram_cell_6t_3 inst_cell_25_20 ( BL20, BLN20, WL25);
sram_cell_6t_3 inst_cell_25_19 ( BL19, BLN19, WL25);
sram_cell_6t_3 inst_cell_25_18 ( BL18, BLN18, WL25);
sram_cell_6t_3 inst_cell_25_17 ( BL17, BLN17, WL25);
sram_cell_6t_3 inst_cell_25_16 ( BL16, BLN16, WL25);
sram_cell_6t_3 inst_cell_25_15 ( BL15, BLN15, WL25);
sram_cell_6t_3 inst_cell_25_14 ( BL14, BLN14, WL25);
sram_cell_6t_3 inst_cell_25_13 ( BL13, BLN13, WL25);
sram_cell_6t_3 inst_cell_25_12 ( BL12, BLN12, WL25);
sram_cell_6t_3 inst_cell_25_11 ( BL11, BLN11, WL25);
sram_cell_6t_3 inst_cell_25_10 ( BL10, BLN10, WL25);
sram_cell_6t_3 inst_cell_25_9 ( BL9, BLN9, WL25);
sram_cell_6t_3 inst_cell_25_8 ( BL8, BLN8, WL25);
sram_cell_6t_3 inst_cell_25_7 ( BL7, BLN7, WL25);
sram_cell_6t_3 inst_cell_25_6 ( BL6, BLN6, WL25);
sram_cell_6t_3 inst_cell_25_5 ( BL5, BLN5, WL25);
sram_cell_6t_3 inst_cell_25_4 ( BL4, BLN4, WL25);
sram_cell_6t_3 inst_cell_25_3 ( BL3, BLN3, WL25);
sram_cell_6t_3 inst_cell_25_2 ( BL2, BLN2, WL25);
sram_cell_6t_3 inst_cell_25_1 ( BL1, BLN1, WL25);
sram_cell_6t_3 inst_cell_25_0 ( BL0, BLN0, WL25);
sram_cell_6t_3 inst_cell_24_127 ( BL127, BLN127, WL24);
sram_cell_6t_3 inst_cell_24_126 ( BL126, BLN126, WL24);
sram_cell_6t_3 inst_cell_24_125 ( BL125, BLN125, WL24);
sram_cell_6t_3 inst_cell_24_124 ( BL124, BLN124, WL24);
sram_cell_6t_3 inst_cell_24_123 ( BL123, BLN123, WL24);
sram_cell_6t_3 inst_cell_24_122 ( BL122, BLN122, WL24);
sram_cell_6t_3 inst_cell_24_121 ( BL121, BLN121, WL24);
sram_cell_6t_3 inst_cell_24_120 ( BL120, BLN120, WL24);
sram_cell_6t_3 inst_cell_24_119 ( BL119, BLN119, WL24);
sram_cell_6t_3 inst_cell_24_118 ( BL118, BLN118, WL24);
sram_cell_6t_3 inst_cell_24_117 ( BL117, BLN117, WL24);
sram_cell_6t_3 inst_cell_24_116 ( BL116, BLN116, WL24);
sram_cell_6t_3 inst_cell_24_115 ( BL115, BLN115, WL24);
sram_cell_6t_3 inst_cell_24_114 ( BL114, BLN114, WL24);
sram_cell_6t_3 inst_cell_24_113 ( BL113, BLN113, WL24);
sram_cell_6t_3 inst_cell_24_112 ( BL112, BLN112, WL24);
sram_cell_6t_3 inst_cell_24_111 ( BL111, BLN111, WL24);
sram_cell_6t_3 inst_cell_24_110 ( BL110, BLN110, WL24);
sram_cell_6t_3 inst_cell_24_109 ( BL109, BLN109, WL24);
sram_cell_6t_3 inst_cell_24_108 ( BL108, BLN108, WL24);
sram_cell_6t_3 inst_cell_24_107 ( BL107, BLN107, WL24);
sram_cell_6t_3 inst_cell_24_106 ( BL106, BLN106, WL24);
sram_cell_6t_3 inst_cell_24_105 ( BL105, BLN105, WL24);
sram_cell_6t_3 inst_cell_24_104 ( BL104, BLN104, WL24);
sram_cell_6t_3 inst_cell_24_103 ( BL103, BLN103, WL24);
sram_cell_6t_3 inst_cell_24_102 ( BL102, BLN102, WL24);
sram_cell_6t_3 inst_cell_24_101 ( BL101, BLN101, WL24);
sram_cell_6t_3 inst_cell_24_100 ( BL100, BLN100, WL24);
sram_cell_6t_3 inst_cell_24_99 ( BL99, BLN99, WL24);
sram_cell_6t_3 inst_cell_24_98 ( BL98, BLN98, WL24);
sram_cell_6t_3 inst_cell_24_97 ( BL97, BLN97, WL24);
sram_cell_6t_3 inst_cell_24_96 ( BL96, BLN96, WL24);
sram_cell_6t_3 inst_cell_24_95 ( BL95, BLN95, WL24);
sram_cell_6t_3 inst_cell_24_94 ( BL94, BLN94, WL24);
sram_cell_6t_3 inst_cell_24_93 ( BL93, BLN93, WL24);
sram_cell_6t_3 inst_cell_24_92 ( BL92, BLN92, WL24);
sram_cell_6t_3 inst_cell_24_91 ( BL91, BLN91, WL24);
sram_cell_6t_3 inst_cell_24_90 ( BL90, BLN90, WL24);
sram_cell_6t_3 inst_cell_24_89 ( BL89, BLN89, WL24);
sram_cell_6t_3 inst_cell_24_88 ( BL88, BLN88, WL24);
sram_cell_6t_3 inst_cell_24_87 ( BL87, BLN87, WL24);
sram_cell_6t_3 inst_cell_24_86 ( BL86, BLN86, WL24);
sram_cell_6t_3 inst_cell_24_85 ( BL85, BLN85, WL24);
sram_cell_6t_3 inst_cell_24_84 ( BL84, BLN84, WL24);
sram_cell_6t_3 inst_cell_24_83 ( BL83, BLN83, WL24);
sram_cell_6t_3 inst_cell_24_82 ( BL82, BLN82, WL24);
sram_cell_6t_3 inst_cell_24_81 ( BL81, BLN81, WL24);
sram_cell_6t_3 inst_cell_24_80 ( BL80, BLN80, WL24);
sram_cell_6t_3 inst_cell_24_79 ( BL79, BLN79, WL24);
sram_cell_6t_3 inst_cell_24_78 ( BL78, BLN78, WL24);
sram_cell_6t_3 inst_cell_24_77 ( BL77, BLN77, WL24);
sram_cell_6t_3 inst_cell_24_76 ( BL76, BLN76, WL24);
sram_cell_6t_3 inst_cell_24_75 ( BL75, BLN75, WL24);
sram_cell_6t_3 inst_cell_24_74 ( BL74, BLN74, WL24);
sram_cell_6t_3 inst_cell_24_73 ( BL73, BLN73, WL24);
sram_cell_6t_3 inst_cell_24_72 ( BL72, BLN72, WL24);
sram_cell_6t_3 inst_cell_24_71 ( BL71, BLN71, WL24);
sram_cell_6t_3 inst_cell_24_70 ( BL70, BLN70, WL24);
sram_cell_6t_3 inst_cell_24_69 ( BL69, BLN69, WL24);
sram_cell_6t_3 inst_cell_24_68 ( BL68, BLN68, WL24);
sram_cell_6t_3 inst_cell_24_67 ( BL67, BLN67, WL24);
sram_cell_6t_3 inst_cell_24_66 ( BL66, BLN66, WL24);
sram_cell_6t_3 inst_cell_24_65 ( BL65, BLN65, WL24);
sram_cell_6t_3 inst_cell_24_64 ( BL64, BLN64, WL24);
sram_cell_6t_3 inst_cell_24_63 ( BL63, BLN63, WL24);
sram_cell_6t_3 inst_cell_24_62 ( BL62, BLN62, WL24);
sram_cell_6t_3 inst_cell_24_61 ( BL61, BLN61, WL24);
sram_cell_6t_3 inst_cell_24_60 ( BL60, BLN60, WL24);
sram_cell_6t_3 inst_cell_24_59 ( BL59, BLN59, WL24);
sram_cell_6t_3 inst_cell_24_58 ( BL58, BLN58, WL24);
sram_cell_6t_3 inst_cell_24_57 ( BL57, BLN57, WL24);
sram_cell_6t_3 inst_cell_24_56 ( BL56, BLN56, WL24);
sram_cell_6t_3 inst_cell_24_55 ( BL55, BLN55, WL24);
sram_cell_6t_3 inst_cell_24_54 ( BL54, BLN54, WL24);
sram_cell_6t_3 inst_cell_24_53 ( BL53, BLN53, WL24);
sram_cell_6t_3 inst_cell_24_52 ( BL52, BLN52, WL24);
sram_cell_6t_3 inst_cell_24_51 ( BL51, BLN51, WL24);
sram_cell_6t_3 inst_cell_24_50 ( BL50, BLN50, WL24);
sram_cell_6t_3 inst_cell_24_49 ( BL49, BLN49, WL24);
sram_cell_6t_3 inst_cell_24_48 ( BL48, BLN48, WL24);
sram_cell_6t_3 inst_cell_24_47 ( BL47, BLN47, WL24);
sram_cell_6t_3 inst_cell_24_46 ( BL46, BLN46, WL24);
sram_cell_6t_3 inst_cell_24_45 ( BL45, BLN45, WL24);
sram_cell_6t_3 inst_cell_24_44 ( BL44, BLN44, WL24);
sram_cell_6t_3 inst_cell_24_43 ( BL43, BLN43, WL24);
sram_cell_6t_3 inst_cell_24_42 ( BL42, BLN42, WL24);
sram_cell_6t_3 inst_cell_24_41 ( BL41, BLN41, WL24);
sram_cell_6t_3 inst_cell_24_40 ( BL40, BLN40, WL24);
sram_cell_6t_3 inst_cell_24_39 ( BL39, BLN39, WL24);
sram_cell_6t_3 inst_cell_24_38 ( BL38, BLN38, WL24);
sram_cell_6t_3 inst_cell_24_37 ( BL37, BLN37, WL24);
sram_cell_6t_3 inst_cell_24_36 ( BL36, BLN36, WL24);
sram_cell_6t_3 inst_cell_24_35 ( BL35, BLN35, WL24);
sram_cell_6t_3 inst_cell_24_34 ( BL34, BLN34, WL24);
sram_cell_6t_3 inst_cell_24_33 ( BL33, BLN33, WL24);
sram_cell_6t_3 inst_cell_24_32 ( BL32, BLN32, WL24);
sram_cell_6t_3 inst_cell_24_31 ( BL31, BLN31, WL24);
sram_cell_6t_3 inst_cell_24_30 ( BL30, BLN30, WL24);
sram_cell_6t_3 inst_cell_24_29 ( BL29, BLN29, WL24);
sram_cell_6t_3 inst_cell_24_28 ( BL28, BLN28, WL24);
sram_cell_6t_3 inst_cell_24_27 ( BL27, BLN27, WL24);
sram_cell_6t_3 inst_cell_24_26 ( BL26, BLN26, WL24);
sram_cell_6t_3 inst_cell_24_25 ( BL25, BLN25, WL24);
sram_cell_6t_3 inst_cell_24_24 ( BL24, BLN24, WL24);
sram_cell_6t_3 inst_cell_24_23 ( BL23, BLN23, WL24);
sram_cell_6t_3 inst_cell_24_22 ( BL22, BLN22, WL24);
sram_cell_6t_3 inst_cell_24_21 ( BL21, BLN21, WL24);
sram_cell_6t_3 inst_cell_24_20 ( BL20, BLN20, WL24);
sram_cell_6t_3 inst_cell_24_19 ( BL19, BLN19, WL24);
sram_cell_6t_3 inst_cell_24_18 ( BL18, BLN18, WL24);
sram_cell_6t_3 inst_cell_24_17 ( BL17, BLN17, WL24);
sram_cell_6t_3 inst_cell_24_16 ( BL16, BLN16, WL24);
sram_cell_6t_3 inst_cell_24_15 ( BL15, BLN15, WL24);
sram_cell_6t_3 inst_cell_24_14 ( BL14, BLN14, WL24);
sram_cell_6t_3 inst_cell_24_13 ( BL13, BLN13, WL24);
sram_cell_6t_3 inst_cell_24_12 ( BL12, BLN12, WL24);
sram_cell_6t_3 inst_cell_24_11 ( BL11, BLN11, WL24);
sram_cell_6t_3 inst_cell_24_10 ( BL10, BLN10, WL24);
sram_cell_6t_3 inst_cell_24_9 ( BL9, BLN9, WL24);
sram_cell_6t_3 inst_cell_24_8 ( BL8, BLN8, WL24);
sram_cell_6t_3 inst_cell_24_7 ( BL7, BLN7, WL24);
sram_cell_6t_3 inst_cell_24_6 ( BL6, BLN6, WL24);
sram_cell_6t_3 inst_cell_24_5 ( BL5, BLN5, WL24);
sram_cell_6t_3 inst_cell_24_4 ( BL4, BLN4, WL24);
sram_cell_6t_3 inst_cell_24_3 ( BL3, BLN3, WL24);
sram_cell_6t_3 inst_cell_24_2 ( BL2, BLN2, WL24);
sram_cell_6t_3 inst_cell_24_1 ( BL1, BLN1, WL24);
sram_cell_6t_3 inst_cell_24_0 ( BL0, BLN0, WL24);
sram_cell_6t_3 inst_cell_23_127 ( BL127, BLN127, WL23);
sram_cell_6t_3 inst_cell_23_126 ( BL126, BLN126, WL23);
sram_cell_6t_3 inst_cell_23_125 ( BL125, BLN125, WL23);
sram_cell_6t_3 inst_cell_23_124 ( BL124, BLN124, WL23);
sram_cell_6t_3 inst_cell_23_123 ( BL123, BLN123, WL23);
sram_cell_6t_3 inst_cell_23_122 ( BL122, BLN122, WL23);
sram_cell_6t_3 inst_cell_23_121 ( BL121, BLN121, WL23);
sram_cell_6t_3 inst_cell_23_120 ( BL120, BLN120, WL23);
sram_cell_6t_3 inst_cell_23_119 ( BL119, BLN119, WL23);
sram_cell_6t_3 inst_cell_23_118 ( BL118, BLN118, WL23);
sram_cell_6t_3 inst_cell_23_117 ( BL117, BLN117, WL23);
sram_cell_6t_3 inst_cell_23_116 ( BL116, BLN116, WL23);
sram_cell_6t_3 inst_cell_23_115 ( BL115, BLN115, WL23);
sram_cell_6t_3 inst_cell_23_114 ( BL114, BLN114, WL23);
sram_cell_6t_3 inst_cell_23_113 ( BL113, BLN113, WL23);
sram_cell_6t_3 inst_cell_23_112 ( BL112, BLN112, WL23);
sram_cell_6t_3 inst_cell_23_111 ( BL111, BLN111, WL23);
sram_cell_6t_3 inst_cell_23_110 ( BL110, BLN110, WL23);
sram_cell_6t_3 inst_cell_23_109 ( BL109, BLN109, WL23);
sram_cell_6t_3 inst_cell_23_108 ( BL108, BLN108, WL23);
sram_cell_6t_3 inst_cell_23_107 ( BL107, BLN107, WL23);
sram_cell_6t_3 inst_cell_23_106 ( BL106, BLN106, WL23);
sram_cell_6t_3 inst_cell_23_105 ( BL105, BLN105, WL23);
sram_cell_6t_3 inst_cell_23_104 ( BL104, BLN104, WL23);
sram_cell_6t_3 inst_cell_23_103 ( BL103, BLN103, WL23);
sram_cell_6t_3 inst_cell_23_102 ( BL102, BLN102, WL23);
sram_cell_6t_3 inst_cell_23_101 ( BL101, BLN101, WL23);
sram_cell_6t_3 inst_cell_23_100 ( BL100, BLN100, WL23);
sram_cell_6t_3 inst_cell_23_99 ( BL99, BLN99, WL23);
sram_cell_6t_3 inst_cell_23_98 ( BL98, BLN98, WL23);
sram_cell_6t_3 inst_cell_23_97 ( BL97, BLN97, WL23);
sram_cell_6t_3 inst_cell_23_96 ( BL96, BLN96, WL23);
sram_cell_6t_3 inst_cell_23_95 ( BL95, BLN95, WL23);
sram_cell_6t_3 inst_cell_23_94 ( BL94, BLN94, WL23);
sram_cell_6t_3 inst_cell_23_93 ( BL93, BLN93, WL23);
sram_cell_6t_3 inst_cell_23_92 ( BL92, BLN92, WL23);
sram_cell_6t_3 inst_cell_23_91 ( BL91, BLN91, WL23);
sram_cell_6t_3 inst_cell_23_90 ( BL90, BLN90, WL23);
sram_cell_6t_3 inst_cell_23_89 ( BL89, BLN89, WL23);
sram_cell_6t_3 inst_cell_23_88 ( BL88, BLN88, WL23);
sram_cell_6t_3 inst_cell_23_87 ( BL87, BLN87, WL23);
sram_cell_6t_3 inst_cell_23_86 ( BL86, BLN86, WL23);
sram_cell_6t_3 inst_cell_23_85 ( BL85, BLN85, WL23);
sram_cell_6t_3 inst_cell_23_84 ( BL84, BLN84, WL23);
sram_cell_6t_3 inst_cell_23_83 ( BL83, BLN83, WL23);
sram_cell_6t_3 inst_cell_23_82 ( BL82, BLN82, WL23);
sram_cell_6t_3 inst_cell_23_81 ( BL81, BLN81, WL23);
sram_cell_6t_3 inst_cell_23_80 ( BL80, BLN80, WL23);
sram_cell_6t_3 inst_cell_23_79 ( BL79, BLN79, WL23);
sram_cell_6t_3 inst_cell_23_78 ( BL78, BLN78, WL23);
sram_cell_6t_3 inst_cell_23_77 ( BL77, BLN77, WL23);
sram_cell_6t_3 inst_cell_23_76 ( BL76, BLN76, WL23);
sram_cell_6t_3 inst_cell_23_75 ( BL75, BLN75, WL23);
sram_cell_6t_3 inst_cell_23_74 ( BL74, BLN74, WL23);
sram_cell_6t_3 inst_cell_23_73 ( BL73, BLN73, WL23);
sram_cell_6t_3 inst_cell_23_72 ( BL72, BLN72, WL23);
sram_cell_6t_3 inst_cell_23_71 ( BL71, BLN71, WL23);
sram_cell_6t_3 inst_cell_23_70 ( BL70, BLN70, WL23);
sram_cell_6t_3 inst_cell_23_69 ( BL69, BLN69, WL23);
sram_cell_6t_3 inst_cell_23_68 ( BL68, BLN68, WL23);
sram_cell_6t_3 inst_cell_23_67 ( BL67, BLN67, WL23);
sram_cell_6t_3 inst_cell_23_66 ( BL66, BLN66, WL23);
sram_cell_6t_3 inst_cell_23_65 ( BL65, BLN65, WL23);
sram_cell_6t_3 inst_cell_23_64 ( BL64, BLN64, WL23);
sram_cell_6t_3 inst_cell_23_63 ( BL63, BLN63, WL23);
sram_cell_6t_3 inst_cell_23_62 ( BL62, BLN62, WL23);
sram_cell_6t_3 inst_cell_23_61 ( BL61, BLN61, WL23);
sram_cell_6t_3 inst_cell_23_60 ( BL60, BLN60, WL23);
sram_cell_6t_3 inst_cell_23_59 ( BL59, BLN59, WL23);
sram_cell_6t_3 inst_cell_23_58 ( BL58, BLN58, WL23);
sram_cell_6t_3 inst_cell_23_57 ( BL57, BLN57, WL23);
sram_cell_6t_3 inst_cell_23_56 ( BL56, BLN56, WL23);
sram_cell_6t_3 inst_cell_23_55 ( BL55, BLN55, WL23);
sram_cell_6t_3 inst_cell_23_54 ( BL54, BLN54, WL23);
sram_cell_6t_3 inst_cell_23_53 ( BL53, BLN53, WL23);
sram_cell_6t_3 inst_cell_23_52 ( BL52, BLN52, WL23);
sram_cell_6t_3 inst_cell_23_51 ( BL51, BLN51, WL23);
sram_cell_6t_3 inst_cell_23_50 ( BL50, BLN50, WL23);
sram_cell_6t_3 inst_cell_23_49 ( BL49, BLN49, WL23);
sram_cell_6t_3 inst_cell_23_48 ( BL48, BLN48, WL23);
sram_cell_6t_3 inst_cell_23_47 ( BL47, BLN47, WL23);
sram_cell_6t_3 inst_cell_23_46 ( BL46, BLN46, WL23);
sram_cell_6t_3 inst_cell_23_45 ( BL45, BLN45, WL23);
sram_cell_6t_3 inst_cell_23_44 ( BL44, BLN44, WL23);
sram_cell_6t_3 inst_cell_23_43 ( BL43, BLN43, WL23);
sram_cell_6t_3 inst_cell_23_42 ( BL42, BLN42, WL23);
sram_cell_6t_3 inst_cell_23_41 ( BL41, BLN41, WL23);
sram_cell_6t_3 inst_cell_23_40 ( BL40, BLN40, WL23);
sram_cell_6t_3 inst_cell_23_39 ( BL39, BLN39, WL23);
sram_cell_6t_3 inst_cell_23_38 ( BL38, BLN38, WL23);
sram_cell_6t_3 inst_cell_23_37 ( BL37, BLN37, WL23);
sram_cell_6t_3 inst_cell_23_36 ( BL36, BLN36, WL23);
sram_cell_6t_3 inst_cell_23_35 ( BL35, BLN35, WL23);
sram_cell_6t_3 inst_cell_23_34 ( BL34, BLN34, WL23);
sram_cell_6t_3 inst_cell_23_33 ( BL33, BLN33, WL23);
sram_cell_6t_3 inst_cell_23_32 ( BL32, BLN32, WL23);
sram_cell_6t_3 inst_cell_23_31 ( BL31, BLN31, WL23);
sram_cell_6t_3 inst_cell_23_30 ( BL30, BLN30, WL23);
sram_cell_6t_3 inst_cell_23_29 ( BL29, BLN29, WL23);
sram_cell_6t_3 inst_cell_23_28 ( BL28, BLN28, WL23);
sram_cell_6t_3 inst_cell_23_27 ( BL27, BLN27, WL23);
sram_cell_6t_3 inst_cell_23_26 ( BL26, BLN26, WL23);
sram_cell_6t_3 inst_cell_23_25 ( BL25, BLN25, WL23);
sram_cell_6t_3 inst_cell_23_24 ( BL24, BLN24, WL23);
sram_cell_6t_3 inst_cell_23_23 ( BL23, BLN23, WL23);
sram_cell_6t_3 inst_cell_23_22 ( BL22, BLN22, WL23);
sram_cell_6t_3 inst_cell_23_21 ( BL21, BLN21, WL23);
sram_cell_6t_3 inst_cell_23_20 ( BL20, BLN20, WL23);
sram_cell_6t_3 inst_cell_23_19 ( BL19, BLN19, WL23);
sram_cell_6t_3 inst_cell_23_18 ( BL18, BLN18, WL23);
sram_cell_6t_3 inst_cell_23_17 ( BL17, BLN17, WL23);
sram_cell_6t_3 inst_cell_23_16 ( BL16, BLN16, WL23);
sram_cell_6t_3 inst_cell_23_15 ( BL15, BLN15, WL23);
sram_cell_6t_3 inst_cell_23_14 ( BL14, BLN14, WL23);
sram_cell_6t_3 inst_cell_23_13 ( BL13, BLN13, WL23);
sram_cell_6t_3 inst_cell_23_12 ( BL12, BLN12, WL23);
sram_cell_6t_3 inst_cell_23_11 ( BL11, BLN11, WL23);
sram_cell_6t_3 inst_cell_23_10 ( BL10, BLN10, WL23);
sram_cell_6t_3 inst_cell_23_9 ( BL9, BLN9, WL23);
sram_cell_6t_3 inst_cell_23_8 ( BL8, BLN8, WL23);
sram_cell_6t_3 inst_cell_23_7 ( BL7, BLN7, WL23);
sram_cell_6t_3 inst_cell_23_6 ( BL6, BLN6, WL23);
sram_cell_6t_3 inst_cell_23_5 ( BL5, BLN5, WL23);
sram_cell_6t_3 inst_cell_23_4 ( BL4, BLN4, WL23);
sram_cell_6t_3 inst_cell_23_3 ( BL3, BLN3, WL23);
sram_cell_6t_3 inst_cell_23_2 ( BL2, BLN2, WL23);
sram_cell_6t_3 inst_cell_23_1 ( BL1, BLN1, WL23);
sram_cell_6t_3 inst_cell_23_0 ( BL0, BLN0, WL23);
sram_cell_6t_3 inst_cell_22_127 ( BL127, BLN127, WL22);
sram_cell_6t_3 inst_cell_22_126 ( BL126, BLN126, WL22);
sram_cell_6t_3 inst_cell_22_125 ( BL125, BLN125, WL22);
sram_cell_6t_3 inst_cell_22_124 ( BL124, BLN124, WL22);
sram_cell_6t_3 inst_cell_22_123 ( BL123, BLN123, WL22);
sram_cell_6t_3 inst_cell_22_122 ( BL122, BLN122, WL22);
sram_cell_6t_3 inst_cell_22_121 ( BL121, BLN121, WL22);
sram_cell_6t_3 inst_cell_22_120 ( BL120, BLN120, WL22);
sram_cell_6t_3 inst_cell_22_119 ( BL119, BLN119, WL22);
sram_cell_6t_3 inst_cell_22_118 ( BL118, BLN118, WL22);
sram_cell_6t_3 inst_cell_22_117 ( BL117, BLN117, WL22);
sram_cell_6t_3 inst_cell_22_116 ( BL116, BLN116, WL22);
sram_cell_6t_3 inst_cell_22_115 ( BL115, BLN115, WL22);
sram_cell_6t_3 inst_cell_22_114 ( BL114, BLN114, WL22);
sram_cell_6t_3 inst_cell_22_113 ( BL113, BLN113, WL22);
sram_cell_6t_3 inst_cell_22_112 ( BL112, BLN112, WL22);
sram_cell_6t_3 inst_cell_22_111 ( BL111, BLN111, WL22);
sram_cell_6t_3 inst_cell_22_110 ( BL110, BLN110, WL22);
sram_cell_6t_3 inst_cell_22_109 ( BL109, BLN109, WL22);
sram_cell_6t_3 inst_cell_22_108 ( BL108, BLN108, WL22);
sram_cell_6t_3 inst_cell_22_107 ( BL107, BLN107, WL22);
sram_cell_6t_3 inst_cell_22_106 ( BL106, BLN106, WL22);
sram_cell_6t_3 inst_cell_22_105 ( BL105, BLN105, WL22);
sram_cell_6t_3 inst_cell_22_104 ( BL104, BLN104, WL22);
sram_cell_6t_3 inst_cell_22_103 ( BL103, BLN103, WL22);
sram_cell_6t_3 inst_cell_22_102 ( BL102, BLN102, WL22);
sram_cell_6t_3 inst_cell_22_101 ( BL101, BLN101, WL22);
sram_cell_6t_3 inst_cell_22_100 ( BL100, BLN100, WL22);
sram_cell_6t_3 inst_cell_22_99 ( BL99, BLN99, WL22);
sram_cell_6t_3 inst_cell_22_98 ( BL98, BLN98, WL22);
sram_cell_6t_3 inst_cell_22_97 ( BL97, BLN97, WL22);
sram_cell_6t_3 inst_cell_22_96 ( BL96, BLN96, WL22);
sram_cell_6t_3 inst_cell_22_95 ( BL95, BLN95, WL22);
sram_cell_6t_3 inst_cell_22_94 ( BL94, BLN94, WL22);
sram_cell_6t_3 inst_cell_22_93 ( BL93, BLN93, WL22);
sram_cell_6t_3 inst_cell_22_92 ( BL92, BLN92, WL22);
sram_cell_6t_3 inst_cell_22_91 ( BL91, BLN91, WL22);
sram_cell_6t_3 inst_cell_22_90 ( BL90, BLN90, WL22);
sram_cell_6t_3 inst_cell_22_89 ( BL89, BLN89, WL22);
sram_cell_6t_3 inst_cell_22_88 ( BL88, BLN88, WL22);
sram_cell_6t_3 inst_cell_22_87 ( BL87, BLN87, WL22);
sram_cell_6t_3 inst_cell_22_86 ( BL86, BLN86, WL22);
sram_cell_6t_3 inst_cell_22_85 ( BL85, BLN85, WL22);
sram_cell_6t_3 inst_cell_22_84 ( BL84, BLN84, WL22);
sram_cell_6t_3 inst_cell_22_83 ( BL83, BLN83, WL22);
sram_cell_6t_3 inst_cell_22_82 ( BL82, BLN82, WL22);
sram_cell_6t_3 inst_cell_22_81 ( BL81, BLN81, WL22);
sram_cell_6t_3 inst_cell_22_80 ( BL80, BLN80, WL22);
sram_cell_6t_3 inst_cell_22_79 ( BL79, BLN79, WL22);
sram_cell_6t_3 inst_cell_22_78 ( BL78, BLN78, WL22);
sram_cell_6t_3 inst_cell_22_77 ( BL77, BLN77, WL22);
sram_cell_6t_3 inst_cell_22_76 ( BL76, BLN76, WL22);
sram_cell_6t_3 inst_cell_22_75 ( BL75, BLN75, WL22);
sram_cell_6t_3 inst_cell_22_74 ( BL74, BLN74, WL22);
sram_cell_6t_3 inst_cell_22_73 ( BL73, BLN73, WL22);
sram_cell_6t_3 inst_cell_22_72 ( BL72, BLN72, WL22);
sram_cell_6t_3 inst_cell_22_71 ( BL71, BLN71, WL22);
sram_cell_6t_3 inst_cell_22_70 ( BL70, BLN70, WL22);
sram_cell_6t_3 inst_cell_22_69 ( BL69, BLN69, WL22);
sram_cell_6t_3 inst_cell_22_68 ( BL68, BLN68, WL22);
sram_cell_6t_3 inst_cell_22_67 ( BL67, BLN67, WL22);
sram_cell_6t_3 inst_cell_22_66 ( BL66, BLN66, WL22);
sram_cell_6t_3 inst_cell_22_65 ( BL65, BLN65, WL22);
sram_cell_6t_3 inst_cell_22_64 ( BL64, BLN64, WL22);
sram_cell_6t_3 inst_cell_22_63 ( BL63, BLN63, WL22);
sram_cell_6t_3 inst_cell_22_62 ( BL62, BLN62, WL22);
sram_cell_6t_3 inst_cell_22_61 ( BL61, BLN61, WL22);
sram_cell_6t_3 inst_cell_22_60 ( BL60, BLN60, WL22);
sram_cell_6t_3 inst_cell_22_59 ( BL59, BLN59, WL22);
sram_cell_6t_3 inst_cell_22_58 ( BL58, BLN58, WL22);
sram_cell_6t_3 inst_cell_22_57 ( BL57, BLN57, WL22);
sram_cell_6t_3 inst_cell_22_56 ( BL56, BLN56, WL22);
sram_cell_6t_3 inst_cell_22_55 ( BL55, BLN55, WL22);
sram_cell_6t_3 inst_cell_22_54 ( BL54, BLN54, WL22);
sram_cell_6t_3 inst_cell_22_53 ( BL53, BLN53, WL22);
sram_cell_6t_3 inst_cell_22_52 ( BL52, BLN52, WL22);
sram_cell_6t_3 inst_cell_22_51 ( BL51, BLN51, WL22);
sram_cell_6t_3 inst_cell_22_50 ( BL50, BLN50, WL22);
sram_cell_6t_3 inst_cell_22_49 ( BL49, BLN49, WL22);
sram_cell_6t_3 inst_cell_22_48 ( BL48, BLN48, WL22);
sram_cell_6t_3 inst_cell_22_47 ( BL47, BLN47, WL22);
sram_cell_6t_3 inst_cell_22_46 ( BL46, BLN46, WL22);
sram_cell_6t_3 inst_cell_22_45 ( BL45, BLN45, WL22);
sram_cell_6t_3 inst_cell_22_44 ( BL44, BLN44, WL22);
sram_cell_6t_3 inst_cell_22_43 ( BL43, BLN43, WL22);
sram_cell_6t_3 inst_cell_22_42 ( BL42, BLN42, WL22);
sram_cell_6t_3 inst_cell_22_41 ( BL41, BLN41, WL22);
sram_cell_6t_3 inst_cell_22_40 ( BL40, BLN40, WL22);
sram_cell_6t_3 inst_cell_22_39 ( BL39, BLN39, WL22);
sram_cell_6t_3 inst_cell_22_38 ( BL38, BLN38, WL22);
sram_cell_6t_3 inst_cell_22_37 ( BL37, BLN37, WL22);
sram_cell_6t_3 inst_cell_22_36 ( BL36, BLN36, WL22);
sram_cell_6t_3 inst_cell_22_35 ( BL35, BLN35, WL22);
sram_cell_6t_3 inst_cell_22_34 ( BL34, BLN34, WL22);
sram_cell_6t_3 inst_cell_22_33 ( BL33, BLN33, WL22);
sram_cell_6t_3 inst_cell_22_32 ( BL32, BLN32, WL22);
sram_cell_6t_3 inst_cell_22_31 ( BL31, BLN31, WL22);
sram_cell_6t_3 inst_cell_22_30 ( BL30, BLN30, WL22);
sram_cell_6t_3 inst_cell_22_29 ( BL29, BLN29, WL22);
sram_cell_6t_3 inst_cell_22_28 ( BL28, BLN28, WL22);
sram_cell_6t_3 inst_cell_22_27 ( BL27, BLN27, WL22);
sram_cell_6t_3 inst_cell_22_26 ( BL26, BLN26, WL22);
sram_cell_6t_3 inst_cell_22_25 ( BL25, BLN25, WL22);
sram_cell_6t_3 inst_cell_22_24 ( BL24, BLN24, WL22);
sram_cell_6t_3 inst_cell_22_23 ( BL23, BLN23, WL22);
sram_cell_6t_3 inst_cell_22_22 ( BL22, BLN22, WL22);
sram_cell_6t_3 inst_cell_22_21 ( BL21, BLN21, WL22);
sram_cell_6t_3 inst_cell_22_20 ( BL20, BLN20, WL22);
sram_cell_6t_3 inst_cell_22_19 ( BL19, BLN19, WL22);
sram_cell_6t_3 inst_cell_22_18 ( BL18, BLN18, WL22);
sram_cell_6t_3 inst_cell_22_17 ( BL17, BLN17, WL22);
sram_cell_6t_3 inst_cell_22_16 ( BL16, BLN16, WL22);
sram_cell_6t_3 inst_cell_22_15 ( BL15, BLN15, WL22);
sram_cell_6t_3 inst_cell_22_14 ( BL14, BLN14, WL22);
sram_cell_6t_3 inst_cell_22_13 ( BL13, BLN13, WL22);
sram_cell_6t_3 inst_cell_22_12 ( BL12, BLN12, WL22);
sram_cell_6t_3 inst_cell_22_11 ( BL11, BLN11, WL22);
sram_cell_6t_3 inst_cell_22_10 ( BL10, BLN10, WL22);
sram_cell_6t_3 inst_cell_22_9 ( BL9, BLN9, WL22);
sram_cell_6t_3 inst_cell_22_8 ( BL8, BLN8, WL22);
sram_cell_6t_3 inst_cell_22_7 ( BL7, BLN7, WL22);
sram_cell_6t_3 inst_cell_22_6 ( BL6, BLN6, WL22);
sram_cell_6t_3 inst_cell_22_5 ( BL5, BLN5, WL22);
sram_cell_6t_3 inst_cell_22_4 ( BL4, BLN4, WL22);
sram_cell_6t_3 inst_cell_22_3 ( BL3, BLN3, WL22);
sram_cell_6t_3 inst_cell_22_2 ( BL2, BLN2, WL22);
sram_cell_6t_3 inst_cell_22_1 ( BL1, BLN1, WL22);
sram_cell_6t_3 inst_cell_22_0 ( BL0, BLN0, WL22);
sram_cell_6t_3 inst_cell_21_127 ( BL127, BLN127, WL21);
sram_cell_6t_3 inst_cell_21_126 ( BL126, BLN126, WL21);
sram_cell_6t_3 inst_cell_21_125 ( BL125, BLN125, WL21);
sram_cell_6t_3 inst_cell_21_124 ( BL124, BLN124, WL21);
sram_cell_6t_3 inst_cell_21_123 ( BL123, BLN123, WL21);
sram_cell_6t_3 inst_cell_21_122 ( BL122, BLN122, WL21);
sram_cell_6t_3 inst_cell_21_121 ( BL121, BLN121, WL21);
sram_cell_6t_3 inst_cell_21_120 ( BL120, BLN120, WL21);
sram_cell_6t_3 inst_cell_21_119 ( BL119, BLN119, WL21);
sram_cell_6t_3 inst_cell_21_118 ( BL118, BLN118, WL21);
sram_cell_6t_3 inst_cell_21_117 ( BL117, BLN117, WL21);
sram_cell_6t_3 inst_cell_21_116 ( BL116, BLN116, WL21);
sram_cell_6t_3 inst_cell_21_115 ( BL115, BLN115, WL21);
sram_cell_6t_3 inst_cell_21_114 ( BL114, BLN114, WL21);
sram_cell_6t_3 inst_cell_21_113 ( BL113, BLN113, WL21);
sram_cell_6t_3 inst_cell_21_112 ( BL112, BLN112, WL21);
sram_cell_6t_3 inst_cell_21_111 ( BL111, BLN111, WL21);
sram_cell_6t_3 inst_cell_21_110 ( BL110, BLN110, WL21);
sram_cell_6t_3 inst_cell_21_109 ( BL109, BLN109, WL21);
sram_cell_6t_3 inst_cell_21_108 ( BL108, BLN108, WL21);
sram_cell_6t_3 inst_cell_21_107 ( BL107, BLN107, WL21);
sram_cell_6t_3 inst_cell_21_106 ( BL106, BLN106, WL21);
sram_cell_6t_3 inst_cell_21_105 ( BL105, BLN105, WL21);
sram_cell_6t_3 inst_cell_21_104 ( BL104, BLN104, WL21);
sram_cell_6t_3 inst_cell_21_103 ( BL103, BLN103, WL21);
sram_cell_6t_3 inst_cell_21_102 ( BL102, BLN102, WL21);
sram_cell_6t_3 inst_cell_21_101 ( BL101, BLN101, WL21);
sram_cell_6t_3 inst_cell_21_100 ( BL100, BLN100, WL21);
sram_cell_6t_3 inst_cell_21_99 ( BL99, BLN99, WL21);
sram_cell_6t_3 inst_cell_21_98 ( BL98, BLN98, WL21);
sram_cell_6t_3 inst_cell_21_97 ( BL97, BLN97, WL21);
sram_cell_6t_3 inst_cell_21_96 ( BL96, BLN96, WL21);
sram_cell_6t_3 inst_cell_21_95 ( BL95, BLN95, WL21);
sram_cell_6t_3 inst_cell_21_94 ( BL94, BLN94, WL21);
sram_cell_6t_3 inst_cell_21_93 ( BL93, BLN93, WL21);
sram_cell_6t_3 inst_cell_21_92 ( BL92, BLN92, WL21);
sram_cell_6t_3 inst_cell_21_91 ( BL91, BLN91, WL21);
sram_cell_6t_3 inst_cell_21_90 ( BL90, BLN90, WL21);
sram_cell_6t_3 inst_cell_21_89 ( BL89, BLN89, WL21);
sram_cell_6t_3 inst_cell_21_88 ( BL88, BLN88, WL21);
sram_cell_6t_3 inst_cell_21_87 ( BL87, BLN87, WL21);
sram_cell_6t_3 inst_cell_21_86 ( BL86, BLN86, WL21);
sram_cell_6t_3 inst_cell_21_85 ( BL85, BLN85, WL21);
sram_cell_6t_3 inst_cell_21_84 ( BL84, BLN84, WL21);
sram_cell_6t_3 inst_cell_21_83 ( BL83, BLN83, WL21);
sram_cell_6t_3 inst_cell_21_82 ( BL82, BLN82, WL21);
sram_cell_6t_3 inst_cell_21_81 ( BL81, BLN81, WL21);
sram_cell_6t_3 inst_cell_21_80 ( BL80, BLN80, WL21);
sram_cell_6t_3 inst_cell_21_79 ( BL79, BLN79, WL21);
sram_cell_6t_3 inst_cell_21_78 ( BL78, BLN78, WL21);
sram_cell_6t_3 inst_cell_21_77 ( BL77, BLN77, WL21);
sram_cell_6t_3 inst_cell_21_76 ( BL76, BLN76, WL21);
sram_cell_6t_3 inst_cell_21_75 ( BL75, BLN75, WL21);
sram_cell_6t_3 inst_cell_21_74 ( BL74, BLN74, WL21);
sram_cell_6t_3 inst_cell_21_73 ( BL73, BLN73, WL21);
sram_cell_6t_3 inst_cell_21_72 ( BL72, BLN72, WL21);
sram_cell_6t_3 inst_cell_21_71 ( BL71, BLN71, WL21);
sram_cell_6t_3 inst_cell_21_70 ( BL70, BLN70, WL21);
sram_cell_6t_3 inst_cell_21_69 ( BL69, BLN69, WL21);
sram_cell_6t_3 inst_cell_21_68 ( BL68, BLN68, WL21);
sram_cell_6t_3 inst_cell_21_67 ( BL67, BLN67, WL21);
sram_cell_6t_3 inst_cell_21_66 ( BL66, BLN66, WL21);
sram_cell_6t_3 inst_cell_21_65 ( BL65, BLN65, WL21);
sram_cell_6t_3 inst_cell_21_64 ( BL64, BLN64, WL21);
sram_cell_6t_3 inst_cell_21_63 ( BL63, BLN63, WL21);
sram_cell_6t_3 inst_cell_21_62 ( BL62, BLN62, WL21);
sram_cell_6t_3 inst_cell_21_61 ( BL61, BLN61, WL21);
sram_cell_6t_3 inst_cell_21_60 ( BL60, BLN60, WL21);
sram_cell_6t_3 inst_cell_21_59 ( BL59, BLN59, WL21);
sram_cell_6t_3 inst_cell_21_58 ( BL58, BLN58, WL21);
sram_cell_6t_3 inst_cell_21_57 ( BL57, BLN57, WL21);
sram_cell_6t_3 inst_cell_21_56 ( BL56, BLN56, WL21);
sram_cell_6t_3 inst_cell_21_55 ( BL55, BLN55, WL21);
sram_cell_6t_3 inst_cell_21_54 ( BL54, BLN54, WL21);
sram_cell_6t_3 inst_cell_21_53 ( BL53, BLN53, WL21);
sram_cell_6t_3 inst_cell_21_52 ( BL52, BLN52, WL21);
sram_cell_6t_3 inst_cell_21_51 ( BL51, BLN51, WL21);
sram_cell_6t_3 inst_cell_21_50 ( BL50, BLN50, WL21);
sram_cell_6t_3 inst_cell_21_49 ( BL49, BLN49, WL21);
sram_cell_6t_3 inst_cell_21_48 ( BL48, BLN48, WL21);
sram_cell_6t_3 inst_cell_21_47 ( BL47, BLN47, WL21);
sram_cell_6t_3 inst_cell_21_46 ( BL46, BLN46, WL21);
sram_cell_6t_3 inst_cell_21_45 ( BL45, BLN45, WL21);
sram_cell_6t_3 inst_cell_21_44 ( BL44, BLN44, WL21);
sram_cell_6t_3 inst_cell_21_43 ( BL43, BLN43, WL21);
sram_cell_6t_3 inst_cell_21_42 ( BL42, BLN42, WL21);
sram_cell_6t_3 inst_cell_21_41 ( BL41, BLN41, WL21);
sram_cell_6t_3 inst_cell_21_40 ( BL40, BLN40, WL21);
sram_cell_6t_3 inst_cell_21_39 ( BL39, BLN39, WL21);
sram_cell_6t_3 inst_cell_21_38 ( BL38, BLN38, WL21);
sram_cell_6t_3 inst_cell_21_37 ( BL37, BLN37, WL21);
sram_cell_6t_3 inst_cell_21_36 ( BL36, BLN36, WL21);
sram_cell_6t_3 inst_cell_21_35 ( BL35, BLN35, WL21);
sram_cell_6t_3 inst_cell_21_34 ( BL34, BLN34, WL21);
sram_cell_6t_3 inst_cell_21_33 ( BL33, BLN33, WL21);
sram_cell_6t_3 inst_cell_21_32 ( BL32, BLN32, WL21);
sram_cell_6t_3 inst_cell_21_31 ( BL31, BLN31, WL21);
sram_cell_6t_3 inst_cell_21_30 ( BL30, BLN30, WL21);
sram_cell_6t_3 inst_cell_21_29 ( BL29, BLN29, WL21);
sram_cell_6t_3 inst_cell_21_28 ( BL28, BLN28, WL21);
sram_cell_6t_3 inst_cell_21_27 ( BL27, BLN27, WL21);
sram_cell_6t_3 inst_cell_21_26 ( BL26, BLN26, WL21);
sram_cell_6t_3 inst_cell_21_25 ( BL25, BLN25, WL21);
sram_cell_6t_3 inst_cell_21_24 ( BL24, BLN24, WL21);
sram_cell_6t_3 inst_cell_21_23 ( BL23, BLN23, WL21);
sram_cell_6t_3 inst_cell_21_22 ( BL22, BLN22, WL21);
sram_cell_6t_3 inst_cell_21_21 ( BL21, BLN21, WL21);
sram_cell_6t_3 inst_cell_21_20 ( BL20, BLN20, WL21);
sram_cell_6t_3 inst_cell_21_19 ( BL19, BLN19, WL21);
sram_cell_6t_3 inst_cell_21_18 ( BL18, BLN18, WL21);
sram_cell_6t_3 inst_cell_21_17 ( BL17, BLN17, WL21);
sram_cell_6t_3 inst_cell_21_16 ( BL16, BLN16, WL21);
sram_cell_6t_3 inst_cell_21_15 ( BL15, BLN15, WL21);
sram_cell_6t_3 inst_cell_21_14 ( BL14, BLN14, WL21);
sram_cell_6t_3 inst_cell_21_13 ( BL13, BLN13, WL21);
sram_cell_6t_3 inst_cell_21_12 ( BL12, BLN12, WL21);
sram_cell_6t_3 inst_cell_21_11 ( BL11, BLN11, WL21);
sram_cell_6t_3 inst_cell_21_10 ( BL10, BLN10, WL21);
sram_cell_6t_3 inst_cell_21_9 ( BL9, BLN9, WL21);
sram_cell_6t_3 inst_cell_21_8 ( BL8, BLN8, WL21);
sram_cell_6t_3 inst_cell_21_7 ( BL7, BLN7, WL21);
sram_cell_6t_3 inst_cell_21_6 ( BL6, BLN6, WL21);
sram_cell_6t_3 inst_cell_21_5 ( BL5, BLN5, WL21);
sram_cell_6t_3 inst_cell_21_4 ( BL4, BLN4, WL21);
sram_cell_6t_3 inst_cell_21_3 ( BL3, BLN3, WL21);
sram_cell_6t_3 inst_cell_21_2 ( BL2, BLN2, WL21);
sram_cell_6t_3 inst_cell_21_1 ( BL1, BLN1, WL21);
sram_cell_6t_3 inst_cell_21_0 ( BL0, BLN0, WL21);
sram_cell_6t_3 inst_cell_20_127 ( BL127, BLN127, WL20);
sram_cell_6t_3 inst_cell_20_126 ( BL126, BLN126, WL20);
sram_cell_6t_3 inst_cell_20_125 ( BL125, BLN125, WL20);
sram_cell_6t_3 inst_cell_20_124 ( BL124, BLN124, WL20);
sram_cell_6t_3 inst_cell_20_123 ( BL123, BLN123, WL20);
sram_cell_6t_3 inst_cell_20_122 ( BL122, BLN122, WL20);
sram_cell_6t_3 inst_cell_20_121 ( BL121, BLN121, WL20);
sram_cell_6t_3 inst_cell_20_120 ( BL120, BLN120, WL20);
sram_cell_6t_3 inst_cell_20_119 ( BL119, BLN119, WL20);
sram_cell_6t_3 inst_cell_20_118 ( BL118, BLN118, WL20);
sram_cell_6t_3 inst_cell_20_117 ( BL117, BLN117, WL20);
sram_cell_6t_3 inst_cell_20_116 ( BL116, BLN116, WL20);
sram_cell_6t_3 inst_cell_20_115 ( BL115, BLN115, WL20);
sram_cell_6t_3 inst_cell_20_114 ( BL114, BLN114, WL20);
sram_cell_6t_3 inst_cell_20_113 ( BL113, BLN113, WL20);
sram_cell_6t_3 inst_cell_20_112 ( BL112, BLN112, WL20);
sram_cell_6t_3 inst_cell_20_111 ( BL111, BLN111, WL20);
sram_cell_6t_3 inst_cell_20_110 ( BL110, BLN110, WL20);
sram_cell_6t_3 inst_cell_20_109 ( BL109, BLN109, WL20);
sram_cell_6t_3 inst_cell_20_108 ( BL108, BLN108, WL20);
sram_cell_6t_3 inst_cell_20_107 ( BL107, BLN107, WL20);
sram_cell_6t_3 inst_cell_20_106 ( BL106, BLN106, WL20);
sram_cell_6t_3 inst_cell_20_105 ( BL105, BLN105, WL20);
sram_cell_6t_3 inst_cell_20_104 ( BL104, BLN104, WL20);
sram_cell_6t_3 inst_cell_20_103 ( BL103, BLN103, WL20);
sram_cell_6t_3 inst_cell_20_102 ( BL102, BLN102, WL20);
sram_cell_6t_3 inst_cell_20_101 ( BL101, BLN101, WL20);
sram_cell_6t_3 inst_cell_20_100 ( BL100, BLN100, WL20);
sram_cell_6t_3 inst_cell_20_99 ( BL99, BLN99, WL20);
sram_cell_6t_3 inst_cell_20_98 ( BL98, BLN98, WL20);
sram_cell_6t_3 inst_cell_20_97 ( BL97, BLN97, WL20);
sram_cell_6t_3 inst_cell_20_96 ( BL96, BLN96, WL20);
sram_cell_6t_3 inst_cell_20_95 ( BL95, BLN95, WL20);
sram_cell_6t_3 inst_cell_20_94 ( BL94, BLN94, WL20);
sram_cell_6t_3 inst_cell_20_93 ( BL93, BLN93, WL20);
sram_cell_6t_3 inst_cell_20_92 ( BL92, BLN92, WL20);
sram_cell_6t_3 inst_cell_20_91 ( BL91, BLN91, WL20);
sram_cell_6t_3 inst_cell_20_90 ( BL90, BLN90, WL20);
sram_cell_6t_3 inst_cell_20_89 ( BL89, BLN89, WL20);
sram_cell_6t_3 inst_cell_20_88 ( BL88, BLN88, WL20);
sram_cell_6t_3 inst_cell_20_87 ( BL87, BLN87, WL20);
sram_cell_6t_3 inst_cell_20_86 ( BL86, BLN86, WL20);
sram_cell_6t_3 inst_cell_20_85 ( BL85, BLN85, WL20);
sram_cell_6t_3 inst_cell_20_84 ( BL84, BLN84, WL20);
sram_cell_6t_3 inst_cell_20_83 ( BL83, BLN83, WL20);
sram_cell_6t_3 inst_cell_20_82 ( BL82, BLN82, WL20);
sram_cell_6t_3 inst_cell_20_81 ( BL81, BLN81, WL20);
sram_cell_6t_3 inst_cell_20_80 ( BL80, BLN80, WL20);
sram_cell_6t_3 inst_cell_20_79 ( BL79, BLN79, WL20);
sram_cell_6t_3 inst_cell_20_78 ( BL78, BLN78, WL20);
sram_cell_6t_3 inst_cell_20_77 ( BL77, BLN77, WL20);
sram_cell_6t_3 inst_cell_20_76 ( BL76, BLN76, WL20);
sram_cell_6t_3 inst_cell_20_75 ( BL75, BLN75, WL20);
sram_cell_6t_3 inst_cell_20_74 ( BL74, BLN74, WL20);
sram_cell_6t_3 inst_cell_20_73 ( BL73, BLN73, WL20);
sram_cell_6t_3 inst_cell_20_72 ( BL72, BLN72, WL20);
sram_cell_6t_3 inst_cell_20_71 ( BL71, BLN71, WL20);
sram_cell_6t_3 inst_cell_20_70 ( BL70, BLN70, WL20);
sram_cell_6t_3 inst_cell_20_69 ( BL69, BLN69, WL20);
sram_cell_6t_3 inst_cell_20_68 ( BL68, BLN68, WL20);
sram_cell_6t_3 inst_cell_20_67 ( BL67, BLN67, WL20);
sram_cell_6t_3 inst_cell_20_66 ( BL66, BLN66, WL20);
sram_cell_6t_3 inst_cell_20_65 ( BL65, BLN65, WL20);
sram_cell_6t_3 inst_cell_20_64 ( BL64, BLN64, WL20);
sram_cell_6t_3 inst_cell_20_63 ( BL63, BLN63, WL20);
sram_cell_6t_3 inst_cell_20_62 ( BL62, BLN62, WL20);
sram_cell_6t_3 inst_cell_20_61 ( BL61, BLN61, WL20);
sram_cell_6t_3 inst_cell_20_60 ( BL60, BLN60, WL20);
sram_cell_6t_3 inst_cell_20_59 ( BL59, BLN59, WL20);
sram_cell_6t_3 inst_cell_20_58 ( BL58, BLN58, WL20);
sram_cell_6t_3 inst_cell_20_57 ( BL57, BLN57, WL20);
sram_cell_6t_3 inst_cell_20_56 ( BL56, BLN56, WL20);
sram_cell_6t_3 inst_cell_20_55 ( BL55, BLN55, WL20);
sram_cell_6t_3 inst_cell_20_54 ( BL54, BLN54, WL20);
sram_cell_6t_3 inst_cell_20_53 ( BL53, BLN53, WL20);
sram_cell_6t_3 inst_cell_20_52 ( BL52, BLN52, WL20);
sram_cell_6t_3 inst_cell_20_51 ( BL51, BLN51, WL20);
sram_cell_6t_3 inst_cell_20_50 ( BL50, BLN50, WL20);
sram_cell_6t_3 inst_cell_20_49 ( BL49, BLN49, WL20);
sram_cell_6t_3 inst_cell_20_48 ( BL48, BLN48, WL20);
sram_cell_6t_3 inst_cell_20_47 ( BL47, BLN47, WL20);
sram_cell_6t_3 inst_cell_20_46 ( BL46, BLN46, WL20);
sram_cell_6t_3 inst_cell_20_45 ( BL45, BLN45, WL20);
sram_cell_6t_3 inst_cell_20_44 ( BL44, BLN44, WL20);
sram_cell_6t_3 inst_cell_20_43 ( BL43, BLN43, WL20);
sram_cell_6t_3 inst_cell_20_42 ( BL42, BLN42, WL20);
sram_cell_6t_3 inst_cell_20_41 ( BL41, BLN41, WL20);
sram_cell_6t_3 inst_cell_20_40 ( BL40, BLN40, WL20);
sram_cell_6t_3 inst_cell_20_39 ( BL39, BLN39, WL20);
sram_cell_6t_3 inst_cell_20_38 ( BL38, BLN38, WL20);
sram_cell_6t_3 inst_cell_20_37 ( BL37, BLN37, WL20);
sram_cell_6t_3 inst_cell_20_36 ( BL36, BLN36, WL20);
sram_cell_6t_3 inst_cell_20_35 ( BL35, BLN35, WL20);
sram_cell_6t_3 inst_cell_20_34 ( BL34, BLN34, WL20);
sram_cell_6t_3 inst_cell_20_33 ( BL33, BLN33, WL20);
sram_cell_6t_3 inst_cell_20_32 ( BL32, BLN32, WL20);
sram_cell_6t_3 inst_cell_20_31 ( BL31, BLN31, WL20);
sram_cell_6t_3 inst_cell_20_30 ( BL30, BLN30, WL20);
sram_cell_6t_3 inst_cell_20_29 ( BL29, BLN29, WL20);
sram_cell_6t_3 inst_cell_20_28 ( BL28, BLN28, WL20);
sram_cell_6t_3 inst_cell_20_27 ( BL27, BLN27, WL20);
sram_cell_6t_3 inst_cell_20_26 ( BL26, BLN26, WL20);
sram_cell_6t_3 inst_cell_20_25 ( BL25, BLN25, WL20);
sram_cell_6t_3 inst_cell_20_24 ( BL24, BLN24, WL20);
sram_cell_6t_3 inst_cell_20_23 ( BL23, BLN23, WL20);
sram_cell_6t_3 inst_cell_20_22 ( BL22, BLN22, WL20);
sram_cell_6t_3 inst_cell_20_21 ( BL21, BLN21, WL20);
sram_cell_6t_3 inst_cell_20_20 ( BL20, BLN20, WL20);
sram_cell_6t_3 inst_cell_20_19 ( BL19, BLN19, WL20);
sram_cell_6t_3 inst_cell_20_18 ( BL18, BLN18, WL20);
sram_cell_6t_3 inst_cell_20_17 ( BL17, BLN17, WL20);
sram_cell_6t_3 inst_cell_20_16 ( BL16, BLN16, WL20);
sram_cell_6t_3 inst_cell_20_15 ( BL15, BLN15, WL20);
sram_cell_6t_3 inst_cell_20_14 ( BL14, BLN14, WL20);
sram_cell_6t_3 inst_cell_20_13 ( BL13, BLN13, WL20);
sram_cell_6t_3 inst_cell_20_12 ( BL12, BLN12, WL20);
sram_cell_6t_3 inst_cell_20_11 ( BL11, BLN11, WL20);
sram_cell_6t_3 inst_cell_20_10 ( BL10, BLN10, WL20);
sram_cell_6t_3 inst_cell_20_9 ( BL9, BLN9, WL20);
sram_cell_6t_3 inst_cell_20_8 ( BL8, BLN8, WL20);
sram_cell_6t_3 inst_cell_20_7 ( BL7, BLN7, WL20);
sram_cell_6t_3 inst_cell_20_6 ( BL6, BLN6, WL20);
sram_cell_6t_3 inst_cell_20_5 ( BL5, BLN5, WL20);
sram_cell_6t_3 inst_cell_20_4 ( BL4, BLN4, WL20);
sram_cell_6t_3 inst_cell_20_3 ( BL3, BLN3, WL20);
sram_cell_6t_3 inst_cell_20_2 ( BL2, BLN2, WL20);
sram_cell_6t_3 inst_cell_20_1 ( BL1, BLN1, WL20);
sram_cell_6t_3 inst_cell_20_0 ( BL0, BLN0, WL20);
sram_cell_6t_3 inst_cell_19_127 ( BL127, BLN127, WL19);
sram_cell_6t_3 inst_cell_19_126 ( BL126, BLN126, WL19);
sram_cell_6t_3 inst_cell_19_125 ( BL125, BLN125, WL19);
sram_cell_6t_3 inst_cell_19_124 ( BL124, BLN124, WL19);
sram_cell_6t_3 inst_cell_19_123 ( BL123, BLN123, WL19);
sram_cell_6t_3 inst_cell_19_122 ( BL122, BLN122, WL19);
sram_cell_6t_3 inst_cell_19_121 ( BL121, BLN121, WL19);
sram_cell_6t_3 inst_cell_19_120 ( BL120, BLN120, WL19);
sram_cell_6t_3 inst_cell_19_119 ( BL119, BLN119, WL19);
sram_cell_6t_3 inst_cell_19_118 ( BL118, BLN118, WL19);
sram_cell_6t_3 inst_cell_19_117 ( BL117, BLN117, WL19);
sram_cell_6t_3 inst_cell_19_116 ( BL116, BLN116, WL19);
sram_cell_6t_3 inst_cell_19_115 ( BL115, BLN115, WL19);
sram_cell_6t_3 inst_cell_19_114 ( BL114, BLN114, WL19);
sram_cell_6t_3 inst_cell_19_113 ( BL113, BLN113, WL19);
sram_cell_6t_3 inst_cell_19_112 ( BL112, BLN112, WL19);
sram_cell_6t_3 inst_cell_19_111 ( BL111, BLN111, WL19);
sram_cell_6t_3 inst_cell_19_110 ( BL110, BLN110, WL19);
sram_cell_6t_3 inst_cell_19_109 ( BL109, BLN109, WL19);
sram_cell_6t_3 inst_cell_19_108 ( BL108, BLN108, WL19);
sram_cell_6t_3 inst_cell_19_107 ( BL107, BLN107, WL19);
sram_cell_6t_3 inst_cell_19_106 ( BL106, BLN106, WL19);
sram_cell_6t_3 inst_cell_19_105 ( BL105, BLN105, WL19);
sram_cell_6t_3 inst_cell_19_104 ( BL104, BLN104, WL19);
sram_cell_6t_3 inst_cell_19_103 ( BL103, BLN103, WL19);
sram_cell_6t_3 inst_cell_19_102 ( BL102, BLN102, WL19);
sram_cell_6t_3 inst_cell_19_101 ( BL101, BLN101, WL19);
sram_cell_6t_3 inst_cell_19_100 ( BL100, BLN100, WL19);
sram_cell_6t_3 inst_cell_19_99 ( BL99, BLN99, WL19);
sram_cell_6t_3 inst_cell_19_98 ( BL98, BLN98, WL19);
sram_cell_6t_3 inst_cell_19_97 ( BL97, BLN97, WL19);
sram_cell_6t_3 inst_cell_19_96 ( BL96, BLN96, WL19);
sram_cell_6t_3 inst_cell_19_95 ( BL95, BLN95, WL19);
sram_cell_6t_3 inst_cell_19_94 ( BL94, BLN94, WL19);
sram_cell_6t_3 inst_cell_19_93 ( BL93, BLN93, WL19);
sram_cell_6t_3 inst_cell_19_92 ( BL92, BLN92, WL19);
sram_cell_6t_3 inst_cell_19_91 ( BL91, BLN91, WL19);
sram_cell_6t_3 inst_cell_19_90 ( BL90, BLN90, WL19);
sram_cell_6t_3 inst_cell_19_89 ( BL89, BLN89, WL19);
sram_cell_6t_3 inst_cell_19_88 ( BL88, BLN88, WL19);
sram_cell_6t_3 inst_cell_19_87 ( BL87, BLN87, WL19);
sram_cell_6t_3 inst_cell_19_86 ( BL86, BLN86, WL19);
sram_cell_6t_3 inst_cell_19_85 ( BL85, BLN85, WL19);
sram_cell_6t_3 inst_cell_19_84 ( BL84, BLN84, WL19);
sram_cell_6t_3 inst_cell_19_83 ( BL83, BLN83, WL19);
sram_cell_6t_3 inst_cell_19_82 ( BL82, BLN82, WL19);
sram_cell_6t_3 inst_cell_19_81 ( BL81, BLN81, WL19);
sram_cell_6t_3 inst_cell_19_80 ( BL80, BLN80, WL19);
sram_cell_6t_3 inst_cell_19_79 ( BL79, BLN79, WL19);
sram_cell_6t_3 inst_cell_19_78 ( BL78, BLN78, WL19);
sram_cell_6t_3 inst_cell_19_77 ( BL77, BLN77, WL19);
sram_cell_6t_3 inst_cell_19_76 ( BL76, BLN76, WL19);
sram_cell_6t_3 inst_cell_19_75 ( BL75, BLN75, WL19);
sram_cell_6t_3 inst_cell_19_74 ( BL74, BLN74, WL19);
sram_cell_6t_3 inst_cell_19_73 ( BL73, BLN73, WL19);
sram_cell_6t_3 inst_cell_19_72 ( BL72, BLN72, WL19);
sram_cell_6t_3 inst_cell_19_71 ( BL71, BLN71, WL19);
sram_cell_6t_3 inst_cell_19_70 ( BL70, BLN70, WL19);
sram_cell_6t_3 inst_cell_19_69 ( BL69, BLN69, WL19);
sram_cell_6t_3 inst_cell_19_68 ( BL68, BLN68, WL19);
sram_cell_6t_3 inst_cell_19_67 ( BL67, BLN67, WL19);
sram_cell_6t_3 inst_cell_19_66 ( BL66, BLN66, WL19);
sram_cell_6t_3 inst_cell_19_65 ( BL65, BLN65, WL19);
sram_cell_6t_3 inst_cell_19_64 ( BL64, BLN64, WL19);
sram_cell_6t_3 inst_cell_19_63 ( BL63, BLN63, WL19);
sram_cell_6t_3 inst_cell_19_62 ( BL62, BLN62, WL19);
sram_cell_6t_3 inst_cell_19_61 ( BL61, BLN61, WL19);
sram_cell_6t_3 inst_cell_19_60 ( BL60, BLN60, WL19);
sram_cell_6t_3 inst_cell_19_59 ( BL59, BLN59, WL19);
sram_cell_6t_3 inst_cell_19_58 ( BL58, BLN58, WL19);
sram_cell_6t_3 inst_cell_19_57 ( BL57, BLN57, WL19);
sram_cell_6t_3 inst_cell_19_56 ( BL56, BLN56, WL19);
sram_cell_6t_3 inst_cell_19_55 ( BL55, BLN55, WL19);
sram_cell_6t_3 inst_cell_19_54 ( BL54, BLN54, WL19);
sram_cell_6t_3 inst_cell_19_53 ( BL53, BLN53, WL19);
sram_cell_6t_3 inst_cell_19_52 ( BL52, BLN52, WL19);
sram_cell_6t_3 inst_cell_19_51 ( BL51, BLN51, WL19);
sram_cell_6t_3 inst_cell_19_50 ( BL50, BLN50, WL19);
sram_cell_6t_3 inst_cell_19_49 ( BL49, BLN49, WL19);
sram_cell_6t_3 inst_cell_19_48 ( BL48, BLN48, WL19);
sram_cell_6t_3 inst_cell_19_47 ( BL47, BLN47, WL19);
sram_cell_6t_3 inst_cell_19_46 ( BL46, BLN46, WL19);
sram_cell_6t_3 inst_cell_19_45 ( BL45, BLN45, WL19);
sram_cell_6t_3 inst_cell_19_44 ( BL44, BLN44, WL19);
sram_cell_6t_3 inst_cell_19_43 ( BL43, BLN43, WL19);
sram_cell_6t_3 inst_cell_19_42 ( BL42, BLN42, WL19);
sram_cell_6t_3 inst_cell_19_41 ( BL41, BLN41, WL19);
sram_cell_6t_3 inst_cell_19_40 ( BL40, BLN40, WL19);
sram_cell_6t_3 inst_cell_19_39 ( BL39, BLN39, WL19);
sram_cell_6t_3 inst_cell_19_38 ( BL38, BLN38, WL19);
sram_cell_6t_3 inst_cell_19_37 ( BL37, BLN37, WL19);
sram_cell_6t_3 inst_cell_19_36 ( BL36, BLN36, WL19);
sram_cell_6t_3 inst_cell_19_35 ( BL35, BLN35, WL19);
sram_cell_6t_3 inst_cell_19_34 ( BL34, BLN34, WL19);
sram_cell_6t_3 inst_cell_19_33 ( BL33, BLN33, WL19);
sram_cell_6t_3 inst_cell_19_32 ( BL32, BLN32, WL19);
sram_cell_6t_3 inst_cell_19_31 ( BL31, BLN31, WL19);
sram_cell_6t_3 inst_cell_19_30 ( BL30, BLN30, WL19);
sram_cell_6t_3 inst_cell_19_29 ( BL29, BLN29, WL19);
sram_cell_6t_3 inst_cell_19_28 ( BL28, BLN28, WL19);
sram_cell_6t_3 inst_cell_19_27 ( BL27, BLN27, WL19);
sram_cell_6t_3 inst_cell_19_26 ( BL26, BLN26, WL19);
sram_cell_6t_3 inst_cell_19_25 ( BL25, BLN25, WL19);
sram_cell_6t_3 inst_cell_19_24 ( BL24, BLN24, WL19);
sram_cell_6t_3 inst_cell_19_23 ( BL23, BLN23, WL19);
sram_cell_6t_3 inst_cell_19_22 ( BL22, BLN22, WL19);
sram_cell_6t_3 inst_cell_19_21 ( BL21, BLN21, WL19);
sram_cell_6t_3 inst_cell_19_20 ( BL20, BLN20, WL19);
sram_cell_6t_3 inst_cell_19_19 ( BL19, BLN19, WL19);
sram_cell_6t_3 inst_cell_19_18 ( BL18, BLN18, WL19);
sram_cell_6t_3 inst_cell_19_17 ( BL17, BLN17, WL19);
sram_cell_6t_3 inst_cell_19_16 ( BL16, BLN16, WL19);
sram_cell_6t_3 inst_cell_19_15 ( BL15, BLN15, WL19);
sram_cell_6t_3 inst_cell_19_14 ( BL14, BLN14, WL19);
sram_cell_6t_3 inst_cell_19_13 ( BL13, BLN13, WL19);
sram_cell_6t_3 inst_cell_19_12 ( BL12, BLN12, WL19);
sram_cell_6t_3 inst_cell_19_11 ( BL11, BLN11, WL19);
sram_cell_6t_3 inst_cell_19_10 ( BL10, BLN10, WL19);
sram_cell_6t_3 inst_cell_19_9 ( BL9, BLN9, WL19);
sram_cell_6t_3 inst_cell_19_8 ( BL8, BLN8, WL19);
sram_cell_6t_3 inst_cell_19_7 ( BL7, BLN7, WL19);
sram_cell_6t_3 inst_cell_19_6 ( BL6, BLN6, WL19);
sram_cell_6t_3 inst_cell_19_5 ( BL5, BLN5, WL19);
sram_cell_6t_3 inst_cell_19_4 ( BL4, BLN4, WL19);
sram_cell_6t_3 inst_cell_19_3 ( BL3, BLN3, WL19);
sram_cell_6t_3 inst_cell_19_2 ( BL2, BLN2, WL19);
sram_cell_6t_3 inst_cell_19_1 ( BL1, BLN1, WL19);
sram_cell_6t_3 inst_cell_19_0 ( BL0, BLN0, WL19);
sram_cell_6t_3 inst_cell_18_127 ( BL127, BLN127, WL18);
sram_cell_6t_3 inst_cell_18_126 ( BL126, BLN126, WL18);
sram_cell_6t_3 inst_cell_18_125 ( BL125, BLN125, WL18);
sram_cell_6t_3 inst_cell_18_124 ( BL124, BLN124, WL18);
sram_cell_6t_3 inst_cell_18_123 ( BL123, BLN123, WL18);
sram_cell_6t_3 inst_cell_18_122 ( BL122, BLN122, WL18);
sram_cell_6t_3 inst_cell_18_121 ( BL121, BLN121, WL18);
sram_cell_6t_3 inst_cell_18_120 ( BL120, BLN120, WL18);
sram_cell_6t_3 inst_cell_18_119 ( BL119, BLN119, WL18);
sram_cell_6t_3 inst_cell_18_118 ( BL118, BLN118, WL18);
sram_cell_6t_3 inst_cell_18_117 ( BL117, BLN117, WL18);
sram_cell_6t_3 inst_cell_18_116 ( BL116, BLN116, WL18);
sram_cell_6t_3 inst_cell_18_115 ( BL115, BLN115, WL18);
sram_cell_6t_3 inst_cell_18_114 ( BL114, BLN114, WL18);
sram_cell_6t_3 inst_cell_18_113 ( BL113, BLN113, WL18);
sram_cell_6t_3 inst_cell_18_112 ( BL112, BLN112, WL18);
sram_cell_6t_3 inst_cell_18_111 ( BL111, BLN111, WL18);
sram_cell_6t_3 inst_cell_18_110 ( BL110, BLN110, WL18);
sram_cell_6t_3 inst_cell_18_109 ( BL109, BLN109, WL18);
sram_cell_6t_3 inst_cell_18_108 ( BL108, BLN108, WL18);
sram_cell_6t_3 inst_cell_18_107 ( BL107, BLN107, WL18);
sram_cell_6t_3 inst_cell_18_106 ( BL106, BLN106, WL18);
sram_cell_6t_3 inst_cell_18_105 ( BL105, BLN105, WL18);
sram_cell_6t_3 inst_cell_18_104 ( BL104, BLN104, WL18);
sram_cell_6t_3 inst_cell_18_103 ( BL103, BLN103, WL18);
sram_cell_6t_3 inst_cell_18_102 ( BL102, BLN102, WL18);
sram_cell_6t_3 inst_cell_18_101 ( BL101, BLN101, WL18);
sram_cell_6t_3 inst_cell_18_100 ( BL100, BLN100, WL18);
sram_cell_6t_3 inst_cell_18_99 ( BL99, BLN99, WL18);
sram_cell_6t_3 inst_cell_18_98 ( BL98, BLN98, WL18);
sram_cell_6t_3 inst_cell_18_97 ( BL97, BLN97, WL18);
sram_cell_6t_3 inst_cell_18_96 ( BL96, BLN96, WL18);
sram_cell_6t_3 inst_cell_18_95 ( BL95, BLN95, WL18);
sram_cell_6t_3 inst_cell_18_94 ( BL94, BLN94, WL18);
sram_cell_6t_3 inst_cell_18_93 ( BL93, BLN93, WL18);
sram_cell_6t_3 inst_cell_18_92 ( BL92, BLN92, WL18);
sram_cell_6t_3 inst_cell_18_91 ( BL91, BLN91, WL18);
sram_cell_6t_3 inst_cell_18_90 ( BL90, BLN90, WL18);
sram_cell_6t_3 inst_cell_18_89 ( BL89, BLN89, WL18);
sram_cell_6t_3 inst_cell_18_88 ( BL88, BLN88, WL18);
sram_cell_6t_3 inst_cell_18_87 ( BL87, BLN87, WL18);
sram_cell_6t_3 inst_cell_18_86 ( BL86, BLN86, WL18);
sram_cell_6t_3 inst_cell_18_85 ( BL85, BLN85, WL18);
sram_cell_6t_3 inst_cell_18_84 ( BL84, BLN84, WL18);
sram_cell_6t_3 inst_cell_18_83 ( BL83, BLN83, WL18);
sram_cell_6t_3 inst_cell_18_82 ( BL82, BLN82, WL18);
sram_cell_6t_3 inst_cell_18_81 ( BL81, BLN81, WL18);
sram_cell_6t_3 inst_cell_18_80 ( BL80, BLN80, WL18);
sram_cell_6t_3 inst_cell_18_79 ( BL79, BLN79, WL18);
sram_cell_6t_3 inst_cell_18_78 ( BL78, BLN78, WL18);
sram_cell_6t_3 inst_cell_18_77 ( BL77, BLN77, WL18);
sram_cell_6t_3 inst_cell_18_76 ( BL76, BLN76, WL18);
sram_cell_6t_3 inst_cell_18_75 ( BL75, BLN75, WL18);
sram_cell_6t_3 inst_cell_18_74 ( BL74, BLN74, WL18);
sram_cell_6t_3 inst_cell_18_73 ( BL73, BLN73, WL18);
sram_cell_6t_3 inst_cell_18_72 ( BL72, BLN72, WL18);
sram_cell_6t_3 inst_cell_18_71 ( BL71, BLN71, WL18);
sram_cell_6t_3 inst_cell_18_70 ( BL70, BLN70, WL18);
sram_cell_6t_3 inst_cell_18_69 ( BL69, BLN69, WL18);
sram_cell_6t_3 inst_cell_18_68 ( BL68, BLN68, WL18);
sram_cell_6t_3 inst_cell_18_67 ( BL67, BLN67, WL18);
sram_cell_6t_3 inst_cell_18_66 ( BL66, BLN66, WL18);
sram_cell_6t_3 inst_cell_18_65 ( BL65, BLN65, WL18);
sram_cell_6t_3 inst_cell_18_64 ( BL64, BLN64, WL18);
sram_cell_6t_3 inst_cell_18_63 ( BL63, BLN63, WL18);
sram_cell_6t_3 inst_cell_18_62 ( BL62, BLN62, WL18);
sram_cell_6t_3 inst_cell_18_61 ( BL61, BLN61, WL18);
sram_cell_6t_3 inst_cell_18_60 ( BL60, BLN60, WL18);
sram_cell_6t_3 inst_cell_18_59 ( BL59, BLN59, WL18);
sram_cell_6t_3 inst_cell_18_58 ( BL58, BLN58, WL18);
sram_cell_6t_3 inst_cell_18_57 ( BL57, BLN57, WL18);
sram_cell_6t_3 inst_cell_18_56 ( BL56, BLN56, WL18);
sram_cell_6t_3 inst_cell_18_55 ( BL55, BLN55, WL18);
sram_cell_6t_3 inst_cell_18_54 ( BL54, BLN54, WL18);
sram_cell_6t_3 inst_cell_18_53 ( BL53, BLN53, WL18);
sram_cell_6t_3 inst_cell_18_52 ( BL52, BLN52, WL18);
sram_cell_6t_3 inst_cell_18_51 ( BL51, BLN51, WL18);
sram_cell_6t_3 inst_cell_18_50 ( BL50, BLN50, WL18);
sram_cell_6t_3 inst_cell_18_49 ( BL49, BLN49, WL18);
sram_cell_6t_3 inst_cell_18_48 ( BL48, BLN48, WL18);
sram_cell_6t_3 inst_cell_18_47 ( BL47, BLN47, WL18);
sram_cell_6t_3 inst_cell_18_46 ( BL46, BLN46, WL18);
sram_cell_6t_3 inst_cell_18_45 ( BL45, BLN45, WL18);
sram_cell_6t_3 inst_cell_18_44 ( BL44, BLN44, WL18);
sram_cell_6t_3 inst_cell_18_43 ( BL43, BLN43, WL18);
sram_cell_6t_3 inst_cell_18_42 ( BL42, BLN42, WL18);
sram_cell_6t_3 inst_cell_18_41 ( BL41, BLN41, WL18);
sram_cell_6t_3 inst_cell_18_40 ( BL40, BLN40, WL18);
sram_cell_6t_3 inst_cell_18_39 ( BL39, BLN39, WL18);
sram_cell_6t_3 inst_cell_18_38 ( BL38, BLN38, WL18);
sram_cell_6t_3 inst_cell_18_37 ( BL37, BLN37, WL18);
sram_cell_6t_3 inst_cell_18_36 ( BL36, BLN36, WL18);
sram_cell_6t_3 inst_cell_18_35 ( BL35, BLN35, WL18);
sram_cell_6t_3 inst_cell_18_34 ( BL34, BLN34, WL18);
sram_cell_6t_3 inst_cell_18_33 ( BL33, BLN33, WL18);
sram_cell_6t_3 inst_cell_18_32 ( BL32, BLN32, WL18);
sram_cell_6t_3 inst_cell_18_31 ( BL31, BLN31, WL18);
sram_cell_6t_3 inst_cell_18_30 ( BL30, BLN30, WL18);
sram_cell_6t_3 inst_cell_18_29 ( BL29, BLN29, WL18);
sram_cell_6t_3 inst_cell_18_28 ( BL28, BLN28, WL18);
sram_cell_6t_3 inst_cell_18_27 ( BL27, BLN27, WL18);
sram_cell_6t_3 inst_cell_18_26 ( BL26, BLN26, WL18);
sram_cell_6t_3 inst_cell_18_25 ( BL25, BLN25, WL18);
sram_cell_6t_3 inst_cell_18_24 ( BL24, BLN24, WL18);
sram_cell_6t_3 inst_cell_18_23 ( BL23, BLN23, WL18);
sram_cell_6t_3 inst_cell_18_22 ( BL22, BLN22, WL18);
sram_cell_6t_3 inst_cell_18_21 ( BL21, BLN21, WL18);
sram_cell_6t_3 inst_cell_18_20 ( BL20, BLN20, WL18);
sram_cell_6t_3 inst_cell_18_19 ( BL19, BLN19, WL18);
sram_cell_6t_3 inst_cell_18_18 ( BL18, BLN18, WL18);
sram_cell_6t_3 inst_cell_18_17 ( BL17, BLN17, WL18);
sram_cell_6t_3 inst_cell_18_16 ( BL16, BLN16, WL18);
sram_cell_6t_3 inst_cell_18_15 ( BL15, BLN15, WL18);
sram_cell_6t_3 inst_cell_18_14 ( BL14, BLN14, WL18);
sram_cell_6t_3 inst_cell_18_13 ( BL13, BLN13, WL18);
sram_cell_6t_3 inst_cell_18_12 ( BL12, BLN12, WL18);
sram_cell_6t_3 inst_cell_18_11 ( BL11, BLN11, WL18);
sram_cell_6t_3 inst_cell_18_10 ( BL10, BLN10, WL18);
sram_cell_6t_3 inst_cell_18_9 ( BL9, BLN9, WL18);
sram_cell_6t_3 inst_cell_18_8 ( BL8, BLN8, WL18);
sram_cell_6t_3 inst_cell_18_7 ( BL7, BLN7, WL18);
sram_cell_6t_3 inst_cell_18_6 ( BL6, BLN6, WL18);
sram_cell_6t_3 inst_cell_18_5 ( BL5, BLN5, WL18);
sram_cell_6t_3 inst_cell_18_4 ( BL4, BLN4, WL18);
sram_cell_6t_3 inst_cell_18_3 ( BL3, BLN3, WL18);
sram_cell_6t_3 inst_cell_18_2 ( BL2, BLN2, WL18);
sram_cell_6t_3 inst_cell_18_1 ( BL1, BLN1, WL18);
sram_cell_6t_3 inst_cell_18_0 ( BL0, BLN0, WL18);
sram_cell_6t_3 inst_cell_17_127 ( BL127, BLN127, WL17);
sram_cell_6t_3 inst_cell_17_126 ( BL126, BLN126, WL17);
sram_cell_6t_3 inst_cell_17_125 ( BL125, BLN125, WL17);
sram_cell_6t_3 inst_cell_17_124 ( BL124, BLN124, WL17);
sram_cell_6t_3 inst_cell_17_123 ( BL123, BLN123, WL17);
sram_cell_6t_3 inst_cell_17_122 ( BL122, BLN122, WL17);
sram_cell_6t_3 inst_cell_17_121 ( BL121, BLN121, WL17);
sram_cell_6t_3 inst_cell_17_120 ( BL120, BLN120, WL17);
sram_cell_6t_3 inst_cell_17_119 ( BL119, BLN119, WL17);
sram_cell_6t_3 inst_cell_17_118 ( BL118, BLN118, WL17);
sram_cell_6t_3 inst_cell_17_117 ( BL117, BLN117, WL17);
sram_cell_6t_3 inst_cell_17_116 ( BL116, BLN116, WL17);
sram_cell_6t_3 inst_cell_17_115 ( BL115, BLN115, WL17);
sram_cell_6t_3 inst_cell_17_114 ( BL114, BLN114, WL17);
sram_cell_6t_3 inst_cell_17_113 ( BL113, BLN113, WL17);
sram_cell_6t_3 inst_cell_17_112 ( BL112, BLN112, WL17);
sram_cell_6t_3 inst_cell_17_111 ( BL111, BLN111, WL17);
sram_cell_6t_3 inst_cell_17_110 ( BL110, BLN110, WL17);
sram_cell_6t_3 inst_cell_17_109 ( BL109, BLN109, WL17);
sram_cell_6t_3 inst_cell_17_108 ( BL108, BLN108, WL17);
sram_cell_6t_3 inst_cell_17_107 ( BL107, BLN107, WL17);
sram_cell_6t_3 inst_cell_17_106 ( BL106, BLN106, WL17);
sram_cell_6t_3 inst_cell_17_105 ( BL105, BLN105, WL17);
sram_cell_6t_3 inst_cell_17_104 ( BL104, BLN104, WL17);
sram_cell_6t_3 inst_cell_17_103 ( BL103, BLN103, WL17);
sram_cell_6t_3 inst_cell_17_102 ( BL102, BLN102, WL17);
sram_cell_6t_3 inst_cell_17_101 ( BL101, BLN101, WL17);
sram_cell_6t_3 inst_cell_17_100 ( BL100, BLN100, WL17);
sram_cell_6t_3 inst_cell_17_99 ( BL99, BLN99, WL17);
sram_cell_6t_3 inst_cell_17_98 ( BL98, BLN98, WL17);
sram_cell_6t_3 inst_cell_17_97 ( BL97, BLN97, WL17);
sram_cell_6t_3 inst_cell_17_96 ( BL96, BLN96, WL17);
sram_cell_6t_3 inst_cell_17_95 ( BL95, BLN95, WL17);
sram_cell_6t_3 inst_cell_17_94 ( BL94, BLN94, WL17);
sram_cell_6t_3 inst_cell_17_93 ( BL93, BLN93, WL17);
sram_cell_6t_3 inst_cell_17_92 ( BL92, BLN92, WL17);
sram_cell_6t_3 inst_cell_17_91 ( BL91, BLN91, WL17);
sram_cell_6t_3 inst_cell_17_90 ( BL90, BLN90, WL17);
sram_cell_6t_3 inst_cell_17_89 ( BL89, BLN89, WL17);
sram_cell_6t_3 inst_cell_17_88 ( BL88, BLN88, WL17);
sram_cell_6t_3 inst_cell_17_87 ( BL87, BLN87, WL17);
sram_cell_6t_3 inst_cell_17_86 ( BL86, BLN86, WL17);
sram_cell_6t_3 inst_cell_17_85 ( BL85, BLN85, WL17);
sram_cell_6t_3 inst_cell_17_84 ( BL84, BLN84, WL17);
sram_cell_6t_3 inst_cell_17_83 ( BL83, BLN83, WL17);
sram_cell_6t_3 inst_cell_17_82 ( BL82, BLN82, WL17);
sram_cell_6t_3 inst_cell_17_81 ( BL81, BLN81, WL17);
sram_cell_6t_3 inst_cell_17_80 ( BL80, BLN80, WL17);
sram_cell_6t_3 inst_cell_17_79 ( BL79, BLN79, WL17);
sram_cell_6t_3 inst_cell_17_78 ( BL78, BLN78, WL17);
sram_cell_6t_3 inst_cell_17_77 ( BL77, BLN77, WL17);
sram_cell_6t_3 inst_cell_17_76 ( BL76, BLN76, WL17);
sram_cell_6t_3 inst_cell_17_75 ( BL75, BLN75, WL17);
sram_cell_6t_3 inst_cell_17_74 ( BL74, BLN74, WL17);
sram_cell_6t_3 inst_cell_17_73 ( BL73, BLN73, WL17);
sram_cell_6t_3 inst_cell_17_72 ( BL72, BLN72, WL17);
sram_cell_6t_3 inst_cell_17_71 ( BL71, BLN71, WL17);
sram_cell_6t_3 inst_cell_17_70 ( BL70, BLN70, WL17);
sram_cell_6t_3 inst_cell_17_69 ( BL69, BLN69, WL17);
sram_cell_6t_3 inst_cell_17_68 ( BL68, BLN68, WL17);
sram_cell_6t_3 inst_cell_17_67 ( BL67, BLN67, WL17);
sram_cell_6t_3 inst_cell_17_66 ( BL66, BLN66, WL17);
sram_cell_6t_3 inst_cell_17_65 ( BL65, BLN65, WL17);
sram_cell_6t_3 inst_cell_17_64 ( BL64, BLN64, WL17);
sram_cell_6t_3 inst_cell_17_63 ( BL63, BLN63, WL17);
sram_cell_6t_3 inst_cell_17_62 ( BL62, BLN62, WL17);
sram_cell_6t_3 inst_cell_17_61 ( BL61, BLN61, WL17);
sram_cell_6t_3 inst_cell_17_60 ( BL60, BLN60, WL17);
sram_cell_6t_3 inst_cell_17_59 ( BL59, BLN59, WL17);
sram_cell_6t_3 inst_cell_17_58 ( BL58, BLN58, WL17);
sram_cell_6t_3 inst_cell_17_57 ( BL57, BLN57, WL17);
sram_cell_6t_3 inst_cell_17_56 ( BL56, BLN56, WL17);
sram_cell_6t_3 inst_cell_17_55 ( BL55, BLN55, WL17);
sram_cell_6t_3 inst_cell_17_54 ( BL54, BLN54, WL17);
sram_cell_6t_3 inst_cell_17_53 ( BL53, BLN53, WL17);
sram_cell_6t_3 inst_cell_17_52 ( BL52, BLN52, WL17);
sram_cell_6t_3 inst_cell_17_51 ( BL51, BLN51, WL17);
sram_cell_6t_3 inst_cell_17_50 ( BL50, BLN50, WL17);
sram_cell_6t_3 inst_cell_17_49 ( BL49, BLN49, WL17);
sram_cell_6t_3 inst_cell_17_48 ( BL48, BLN48, WL17);
sram_cell_6t_3 inst_cell_17_47 ( BL47, BLN47, WL17);
sram_cell_6t_3 inst_cell_17_46 ( BL46, BLN46, WL17);
sram_cell_6t_3 inst_cell_17_45 ( BL45, BLN45, WL17);
sram_cell_6t_3 inst_cell_17_44 ( BL44, BLN44, WL17);
sram_cell_6t_3 inst_cell_17_43 ( BL43, BLN43, WL17);
sram_cell_6t_3 inst_cell_17_42 ( BL42, BLN42, WL17);
sram_cell_6t_3 inst_cell_17_41 ( BL41, BLN41, WL17);
sram_cell_6t_3 inst_cell_17_40 ( BL40, BLN40, WL17);
sram_cell_6t_3 inst_cell_17_39 ( BL39, BLN39, WL17);
sram_cell_6t_3 inst_cell_17_38 ( BL38, BLN38, WL17);
sram_cell_6t_3 inst_cell_17_37 ( BL37, BLN37, WL17);
sram_cell_6t_3 inst_cell_17_36 ( BL36, BLN36, WL17);
sram_cell_6t_3 inst_cell_17_35 ( BL35, BLN35, WL17);
sram_cell_6t_3 inst_cell_17_34 ( BL34, BLN34, WL17);
sram_cell_6t_3 inst_cell_17_33 ( BL33, BLN33, WL17);
sram_cell_6t_3 inst_cell_17_32 ( BL32, BLN32, WL17);
sram_cell_6t_3 inst_cell_17_31 ( BL31, BLN31, WL17);
sram_cell_6t_3 inst_cell_17_30 ( BL30, BLN30, WL17);
sram_cell_6t_3 inst_cell_17_29 ( BL29, BLN29, WL17);
sram_cell_6t_3 inst_cell_17_28 ( BL28, BLN28, WL17);
sram_cell_6t_3 inst_cell_17_27 ( BL27, BLN27, WL17);
sram_cell_6t_3 inst_cell_17_26 ( BL26, BLN26, WL17);
sram_cell_6t_3 inst_cell_17_25 ( BL25, BLN25, WL17);
sram_cell_6t_3 inst_cell_17_24 ( BL24, BLN24, WL17);
sram_cell_6t_3 inst_cell_17_23 ( BL23, BLN23, WL17);
sram_cell_6t_3 inst_cell_17_22 ( BL22, BLN22, WL17);
sram_cell_6t_3 inst_cell_17_21 ( BL21, BLN21, WL17);
sram_cell_6t_3 inst_cell_17_20 ( BL20, BLN20, WL17);
sram_cell_6t_3 inst_cell_17_19 ( BL19, BLN19, WL17);
sram_cell_6t_3 inst_cell_17_18 ( BL18, BLN18, WL17);
sram_cell_6t_3 inst_cell_17_17 ( BL17, BLN17, WL17);
sram_cell_6t_3 inst_cell_17_16 ( BL16, BLN16, WL17);
sram_cell_6t_3 inst_cell_17_15 ( BL15, BLN15, WL17);
sram_cell_6t_3 inst_cell_17_14 ( BL14, BLN14, WL17);
sram_cell_6t_3 inst_cell_17_13 ( BL13, BLN13, WL17);
sram_cell_6t_3 inst_cell_17_12 ( BL12, BLN12, WL17);
sram_cell_6t_3 inst_cell_17_11 ( BL11, BLN11, WL17);
sram_cell_6t_3 inst_cell_17_10 ( BL10, BLN10, WL17);
sram_cell_6t_3 inst_cell_17_9 ( BL9, BLN9, WL17);
sram_cell_6t_3 inst_cell_17_8 ( BL8, BLN8, WL17);
sram_cell_6t_3 inst_cell_17_7 ( BL7, BLN7, WL17);
sram_cell_6t_3 inst_cell_17_6 ( BL6, BLN6, WL17);
sram_cell_6t_3 inst_cell_17_5 ( BL5, BLN5, WL17);
sram_cell_6t_3 inst_cell_17_4 ( BL4, BLN4, WL17);
sram_cell_6t_3 inst_cell_17_3 ( BL3, BLN3, WL17);
sram_cell_6t_3 inst_cell_17_2 ( BL2, BLN2, WL17);
sram_cell_6t_3 inst_cell_17_1 ( BL1, BLN1, WL17);
sram_cell_6t_3 inst_cell_17_0 ( BL0, BLN0, WL17);
sram_cell_6t_3 inst_cell_16_127 ( BL127, BLN127, WL16);
sram_cell_6t_3 inst_cell_16_126 ( BL126, BLN126, WL16);
sram_cell_6t_3 inst_cell_16_125 ( BL125, BLN125, WL16);
sram_cell_6t_3 inst_cell_16_124 ( BL124, BLN124, WL16);
sram_cell_6t_3 inst_cell_16_123 ( BL123, BLN123, WL16);
sram_cell_6t_3 inst_cell_16_122 ( BL122, BLN122, WL16);
sram_cell_6t_3 inst_cell_16_121 ( BL121, BLN121, WL16);
sram_cell_6t_3 inst_cell_16_120 ( BL120, BLN120, WL16);
sram_cell_6t_3 inst_cell_16_119 ( BL119, BLN119, WL16);
sram_cell_6t_3 inst_cell_16_118 ( BL118, BLN118, WL16);
sram_cell_6t_3 inst_cell_16_117 ( BL117, BLN117, WL16);
sram_cell_6t_3 inst_cell_16_116 ( BL116, BLN116, WL16);
sram_cell_6t_3 inst_cell_16_115 ( BL115, BLN115, WL16);
sram_cell_6t_3 inst_cell_16_114 ( BL114, BLN114, WL16);
sram_cell_6t_3 inst_cell_16_113 ( BL113, BLN113, WL16);
sram_cell_6t_3 inst_cell_16_112 ( BL112, BLN112, WL16);
sram_cell_6t_3 inst_cell_16_111 ( BL111, BLN111, WL16);
sram_cell_6t_3 inst_cell_16_110 ( BL110, BLN110, WL16);
sram_cell_6t_3 inst_cell_16_109 ( BL109, BLN109, WL16);
sram_cell_6t_3 inst_cell_16_108 ( BL108, BLN108, WL16);
sram_cell_6t_3 inst_cell_16_107 ( BL107, BLN107, WL16);
sram_cell_6t_3 inst_cell_16_106 ( BL106, BLN106, WL16);
sram_cell_6t_3 inst_cell_16_105 ( BL105, BLN105, WL16);
sram_cell_6t_3 inst_cell_16_104 ( BL104, BLN104, WL16);
sram_cell_6t_3 inst_cell_16_103 ( BL103, BLN103, WL16);
sram_cell_6t_3 inst_cell_16_102 ( BL102, BLN102, WL16);
sram_cell_6t_3 inst_cell_16_101 ( BL101, BLN101, WL16);
sram_cell_6t_3 inst_cell_16_100 ( BL100, BLN100, WL16);
sram_cell_6t_3 inst_cell_16_99 ( BL99, BLN99, WL16);
sram_cell_6t_3 inst_cell_16_98 ( BL98, BLN98, WL16);
sram_cell_6t_3 inst_cell_16_97 ( BL97, BLN97, WL16);
sram_cell_6t_3 inst_cell_16_96 ( BL96, BLN96, WL16);
sram_cell_6t_3 inst_cell_16_95 ( BL95, BLN95, WL16);
sram_cell_6t_3 inst_cell_16_94 ( BL94, BLN94, WL16);
sram_cell_6t_3 inst_cell_16_93 ( BL93, BLN93, WL16);
sram_cell_6t_3 inst_cell_16_92 ( BL92, BLN92, WL16);
sram_cell_6t_3 inst_cell_16_91 ( BL91, BLN91, WL16);
sram_cell_6t_3 inst_cell_16_90 ( BL90, BLN90, WL16);
sram_cell_6t_3 inst_cell_16_89 ( BL89, BLN89, WL16);
sram_cell_6t_3 inst_cell_16_88 ( BL88, BLN88, WL16);
sram_cell_6t_3 inst_cell_16_87 ( BL87, BLN87, WL16);
sram_cell_6t_3 inst_cell_16_86 ( BL86, BLN86, WL16);
sram_cell_6t_3 inst_cell_16_85 ( BL85, BLN85, WL16);
sram_cell_6t_3 inst_cell_16_84 ( BL84, BLN84, WL16);
sram_cell_6t_3 inst_cell_16_83 ( BL83, BLN83, WL16);
sram_cell_6t_3 inst_cell_16_82 ( BL82, BLN82, WL16);
sram_cell_6t_3 inst_cell_16_81 ( BL81, BLN81, WL16);
sram_cell_6t_3 inst_cell_16_80 ( BL80, BLN80, WL16);
sram_cell_6t_3 inst_cell_16_79 ( BL79, BLN79, WL16);
sram_cell_6t_3 inst_cell_16_78 ( BL78, BLN78, WL16);
sram_cell_6t_3 inst_cell_16_77 ( BL77, BLN77, WL16);
sram_cell_6t_3 inst_cell_16_76 ( BL76, BLN76, WL16);
sram_cell_6t_3 inst_cell_16_75 ( BL75, BLN75, WL16);
sram_cell_6t_3 inst_cell_16_74 ( BL74, BLN74, WL16);
sram_cell_6t_3 inst_cell_16_73 ( BL73, BLN73, WL16);
sram_cell_6t_3 inst_cell_16_72 ( BL72, BLN72, WL16);
sram_cell_6t_3 inst_cell_16_71 ( BL71, BLN71, WL16);
sram_cell_6t_3 inst_cell_16_70 ( BL70, BLN70, WL16);
sram_cell_6t_3 inst_cell_16_69 ( BL69, BLN69, WL16);
sram_cell_6t_3 inst_cell_16_68 ( BL68, BLN68, WL16);
sram_cell_6t_3 inst_cell_16_67 ( BL67, BLN67, WL16);
sram_cell_6t_3 inst_cell_16_66 ( BL66, BLN66, WL16);
sram_cell_6t_3 inst_cell_16_65 ( BL65, BLN65, WL16);
sram_cell_6t_3 inst_cell_16_64 ( BL64, BLN64, WL16);
sram_cell_6t_3 inst_cell_16_63 ( BL63, BLN63, WL16);
sram_cell_6t_3 inst_cell_16_62 ( BL62, BLN62, WL16);
sram_cell_6t_3 inst_cell_16_61 ( BL61, BLN61, WL16);
sram_cell_6t_3 inst_cell_16_60 ( BL60, BLN60, WL16);
sram_cell_6t_3 inst_cell_16_59 ( BL59, BLN59, WL16);
sram_cell_6t_3 inst_cell_16_58 ( BL58, BLN58, WL16);
sram_cell_6t_3 inst_cell_16_57 ( BL57, BLN57, WL16);
sram_cell_6t_3 inst_cell_16_56 ( BL56, BLN56, WL16);
sram_cell_6t_3 inst_cell_16_55 ( BL55, BLN55, WL16);
sram_cell_6t_3 inst_cell_16_54 ( BL54, BLN54, WL16);
sram_cell_6t_3 inst_cell_16_53 ( BL53, BLN53, WL16);
sram_cell_6t_3 inst_cell_16_52 ( BL52, BLN52, WL16);
sram_cell_6t_3 inst_cell_16_51 ( BL51, BLN51, WL16);
sram_cell_6t_3 inst_cell_16_50 ( BL50, BLN50, WL16);
sram_cell_6t_3 inst_cell_16_49 ( BL49, BLN49, WL16);
sram_cell_6t_3 inst_cell_16_48 ( BL48, BLN48, WL16);
sram_cell_6t_3 inst_cell_16_47 ( BL47, BLN47, WL16);
sram_cell_6t_3 inst_cell_16_46 ( BL46, BLN46, WL16);
sram_cell_6t_3 inst_cell_16_45 ( BL45, BLN45, WL16);
sram_cell_6t_3 inst_cell_16_44 ( BL44, BLN44, WL16);
sram_cell_6t_3 inst_cell_16_43 ( BL43, BLN43, WL16);
sram_cell_6t_3 inst_cell_16_42 ( BL42, BLN42, WL16);
sram_cell_6t_3 inst_cell_16_41 ( BL41, BLN41, WL16);
sram_cell_6t_3 inst_cell_16_40 ( BL40, BLN40, WL16);
sram_cell_6t_3 inst_cell_16_39 ( BL39, BLN39, WL16);
sram_cell_6t_3 inst_cell_16_38 ( BL38, BLN38, WL16);
sram_cell_6t_3 inst_cell_16_37 ( BL37, BLN37, WL16);
sram_cell_6t_3 inst_cell_16_36 ( BL36, BLN36, WL16);
sram_cell_6t_3 inst_cell_16_35 ( BL35, BLN35, WL16);
sram_cell_6t_3 inst_cell_16_34 ( BL34, BLN34, WL16);
sram_cell_6t_3 inst_cell_16_33 ( BL33, BLN33, WL16);
sram_cell_6t_3 inst_cell_16_32 ( BL32, BLN32, WL16);
sram_cell_6t_3 inst_cell_16_31 ( BL31, BLN31, WL16);
sram_cell_6t_3 inst_cell_16_30 ( BL30, BLN30, WL16);
sram_cell_6t_3 inst_cell_16_29 ( BL29, BLN29, WL16);
sram_cell_6t_3 inst_cell_16_28 ( BL28, BLN28, WL16);
sram_cell_6t_3 inst_cell_16_27 ( BL27, BLN27, WL16);
sram_cell_6t_3 inst_cell_16_26 ( BL26, BLN26, WL16);
sram_cell_6t_3 inst_cell_16_25 ( BL25, BLN25, WL16);
sram_cell_6t_3 inst_cell_16_24 ( BL24, BLN24, WL16);
sram_cell_6t_3 inst_cell_16_23 ( BL23, BLN23, WL16);
sram_cell_6t_3 inst_cell_16_22 ( BL22, BLN22, WL16);
sram_cell_6t_3 inst_cell_16_21 ( BL21, BLN21, WL16);
sram_cell_6t_3 inst_cell_16_20 ( BL20, BLN20, WL16);
sram_cell_6t_3 inst_cell_16_19 ( BL19, BLN19, WL16);
sram_cell_6t_3 inst_cell_16_18 ( BL18, BLN18, WL16);
sram_cell_6t_3 inst_cell_16_17 ( BL17, BLN17, WL16);
sram_cell_6t_3 inst_cell_16_16 ( BL16, BLN16, WL16);
sram_cell_6t_3 inst_cell_16_15 ( BL15, BLN15, WL16);
sram_cell_6t_3 inst_cell_16_14 ( BL14, BLN14, WL16);
sram_cell_6t_3 inst_cell_16_13 ( BL13, BLN13, WL16);
sram_cell_6t_3 inst_cell_16_12 ( BL12, BLN12, WL16);
sram_cell_6t_3 inst_cell_16_11 ( BL11, BLN11, WL16);
sram_cell_6t_3 inst_cell_16_10 ( BL10, BLN10, WL16);
sram_cell_6t_3 inst_cell_16_9 ( BL9, BLN9, WL16);
sram_cell_6t_3 inst_cell_16_8 ( BL8, BLN8, WL16);
sram_cell_6t_3 inst_cell_16_7 ( BL7, BLN7, WL16);
sram_cell_6t_3 inst_cell_16_6 ( BL6, BLN6, WL16);
sram_cell_6t_3 inst_cell_16_5 ( BL5, BLN5, WL16);
sram_cell_6t_3 inst_cell_16_4 ( BL4, BLN4, WL16);
sram_cell_6t_3 inst_cell_16_3 ( BL3, BLN3, WL16);
sram_cell_6t_3 inst_cell_16_2 ( BL2, BLN2, WL16);
sram_cell_6t_3 inst_cell_16_1 ( BL1, BLN1, WL16);
sram_cell_6t_3 inst_cell_16_0 ( BL0, BLN0, WL16);
sram_cell_6t_3 inst_cell_15_127 ( BL127, BLN127, WL15);
sram_cell_6t_3 inst_cell_15_126 ( BL126, BLN126, WL15);
sram_cell_6t_3 inst_cell_15_125 ( BL125, BLN125, WL15);
sram_cell_6t_3 inst_cell_15_124 ( BL124, BLN124, WL15);
sram_cell_6t_3 inst_cell_15_123 ( BL123, BLN123, WL15);
sram_cell_6t_3 inst_cell_15_122 ( BL122, BLN122, WL15);
sram_cell_6t_3 inst_cell_15_121 ( BL121, BLN121, WL15);
sram_cell_6t_3 inst_cell_15_120 ( BL120, BLN120, WL15);
sram_cell_6t_3 inst_cell_15_119 ( BL119, BLN119, WL15);
sram_cell_6t_3 inst_cell_15_118 ( BL118, BLN118, WL15);
sram_cell_6t_3 inst_cell_15_117 ( BL117, BLN117, WL15);
sram_cell_6t_3 inst_cell_15_116 ( BL116, BLN116, WL15);
sram_cell_6t_3 inst_cell_15_115 ( BL115, BLN115, WL15);
sram_cell_6t_3 inst_cell_15_114 ( BL114, BLN114, WL15);
sram_cell_6t_3 inst_cell_15_113 ( BL113, BLN113, WL15);
sram_cell_6t_3 inst_cell_15_112 ( BL112, BLN112, WL15);
sram_cell_6t_3 inst_cell_15_111 ( BL111, BLN111, WL15);
sram_cell_6t_3 inst_cell_15_110 ( BL110, BLN110, WL15);
sram_cell_6t_3 inst_cell_15_109 ( BL109, BLN109, WL15);
sram_cell_6t_3 inst_cell_15_108 ( BL108, BLN108, WL15);
sram_cell_6t_3 inst_cell_15_107 ( BL107, BLN107, WL15);
sram_cell_6t_3 inst_cell_15_106 ( BL106, BLN106, WL15);
sram_cell_6t_3 inst_cell_15_105 ( BL105, BLN105, WL15);
sram_cell_6t_3 inst_cell_15_104 ( BL104, BLN104, WL15);
sram_cell_6t_3 inst_cell_15_103 ( BL103, BLN103, WL15);
sram_cell_6t_3 inst_cell_15_102 ( BL102, BLN102, WL15);
sram_cell_6t_3 inst_cell_15_101 ( BL101, BLN101, WL15);
sram_cell_6t_3 inst_cell_15_100 ( BL100, BLN100, WL15);
sram_cell_6t_3 inst_cell_15_99 ( BL99, BLN99, WL15);
sram_cell_6t_3 inst_cell_15_98 ( BL98, BLN98, WL15);
sram_cell_6t_3 inst_cell_15_97 ( BL97, BLN97, WL15);
sram_cell_6t_3 inst_cell_15_96 ( BL96, BLN96, WL15);
sram_cell_6t_3 inst_cell_15_95 ( BL95, BLN95, WL15);
sram_cell_6t_3 inst_cell_15_94 ( BL94, BLN94, WL15);
sram_cell_6t_3 inst_cell_15_93 ( BL93, BLN93, WL15);
sram_cell_6t_3 inst_cell_15_92 ( BL92, BLN92, WL15);
sram_cell_6t_3 inst_cell_15_91 ( BL91, BLN91, WL15);
sram_cell_6t_3 inst_cell_15_90 ( BL90, BLN90, WL15);
sram_cell_6t_3 inst_cell_15_89 ( BL89, BLN89, WL15);
sram_cell_6t_3 inst_cell_15_88 ( BL88, BLN88, WL15);
sram_cell_6t_3 inst_cell_15_87 ( BL87, BLN87, WL15);
sram_cell_6t_3 inst_cell_15_86 ( BL86, BLN86, WL15);
sram_cell_6t_3 inst_cell_15_85 ( BL85, BLN85, WL15);
sram_cell_6t_3 inst_cell_15_84 ( BL84, BLN84, WL15);
sram_cell_6t_3 inst_cell_15_83 ( BL83, BLN83, WL15);
sram_cell_6t_3 inst_cell_15_82 ( BL82, BLN82, WL15);
sram_cell_6t_3 inst_cell_15_81 ( BL81, BLN81, WL15);
sram_cell_6t_3 inst_cell_15_80 ( BL80, BLN80, WL15);
sram_cell_6t_3 inst_cell_15_79 ( BL79, BLN79, WL15);
sram_cell_6t_3 inst_cell_15_78 ( BL78, BLN78, WL15);
sram_cell_6t_3 inst_cell_15_77 ( BL77, BLN77, WL15);
sram_cell_6t_3 inst_cell_15_76 ( BL76, BLN76, WL15);
sram_cell_6t_3 inst_cell_15_75 ( BL75, BLN75, WL15);
sram_cell_6t_3 inst_cell_15_74 ( BL74, BLN74, WL15);
sram_cell_6t_3 inst_cell_15_73 ( BL73, BLN73, WL15);
sram_cell_6t_3 inst_cell_15_72 ( BL72, BLN72, WL15);
sram_cell_6t_3 inst_cell_15_71 ( BL71, BLN71, WL15);
sram_cell_6t_3 inst_cell_15_70 ( BL70, BLN70, WL15);
sram_cell_6t_3 inst_cell_15_69 ( BL69, BLN69, WL15);
sram_cell_6t_3 inst_cell_15_68 ( BL68, BLN68, WL15);
sram_cell_6t_3 inst_cell_15_67 ( BL67, BLN67, WL15);
sram_cell_6t_3 inst_cell_15_66 ( BL66, BLN66, WL15);
sram_cell_6t_3 inst_cell_15_65 ( BL65, BLN65, WL15);
sram_cell_6t_3 inst_cell_15_64 ( BL64, BLN64, WL15);
sram_cell_6t_3 inst_cell_15_63 ( BL63, BLN63, WL15);
sram_cell_6t_3 inst_cell_15_62 ( BL62, BLN62, WL15);
sram_cell_6t_3 inst_cell_15_61 ( BL61, BLN61, WL15);
sram_cell_6t_3 inst_cell_15_60 ( BL60, BLN60, WL15);
sram_cell_6t_3 inst_cell_15_59 ( BL59, BLN59, WL15);
sram_cell_6t_3 inst_cell_15_58 ( BL58, BLN58, WL15);
sram_cell_6t_3 inst_cell_15_57 ( BL57, BLN57, WL15);
sram_cell_6t_3 inst_cell_15_56 ( BL56, BLN56, WL15);
sram_cell_6t_3 inst_cell_15_55 ( BL55, BLN55, WL15);
sram_cell_6t_3 inst_cell_15_54 ( BL54, BLN54, WL15);
sram_cell_6t_3 inst_cell_15_53 ( BL53, BLN53, WL15);
sram_cell_6t_3 inst_cell_15_52 ( BL52, BLN52, WL15);
sram_cell_6t_3 inst_cell_15_51 ( BL51, BLN51, WL15);
sram_cell_6t_3 inst_cell_15_50 ( BL50, BLN50, WL15);
sram_cell_6t_3 inst_cell_15_49 ( BL49, BLN49, WL15);
sram_cell_6t_3 inst_cell_15_48 ( BL48, BLN48, WL15);
sram_cell_6t_3 inst_cell_15_47 ( BL47, BLN47, WL15);
sram_cell_6t_3 inst_cell_15_46 ( BL46, BLN46, WL15);
sram_cell_6t_3 inst_cell_15_45 ( BL45, BLN45, WL15);
sram_cell_6t_3 inst_cell_15_44 ( BL44, BLN44, WL15);
sram_cell_6t_3 inst_cell_15_43 ( BL43, BLN43, WL15);
sram_cell_6t_3 inst_cell_15_42 ( BL42, BLN42, WL15);
sram_cell_6t_3 inst_cell_15_41 ( BL41, BLN41, WL15);
sram_cell_6t_3 inst_cell_15_40 ( BL40, BLN40, WL15);
sram_cell_6t_3 inst_cell_15_39 ( BL39, BLN39, WL15);
sram_cell_6t_3 inst_cell_15_38 ( BL38, BLN38, WL15);
sram_cell_6t_3 inst_cell_15_37 ( BL37, BLN37, WL15);
sram_cell_6t_3 inst_cell_15_36 ( BL36, BLN36, WL15);
sram_cell_6t_3 inst_cell_15_35 ( BL35, BLN35, WL15);
sram_cell_6t_3 inst_cell_15_34 ( BL34, BLN34, WL15);
sram_cell_6t_3 inst_cell_15_33 ( BL33, BLN33, WL15);
sram_cell_6t_3 inst_cell_15_32 ( BL32, BLN32, WL15);
sram_cell_6t_3 inst_cell_15_31 ( BL31, BLN31, WL15);
sram_cell_6t_3 inst_cell_15_30 ( BL30, BLN30, WL15);
sram_cell_6t_3 inst_cell_15_29 ( BL29, BLN29, WL15);
sram_cell_6t_3 inst_cell_15_28 ( BL28, BLN28, WL15);
sram_cell_6t_3 inst_cell_15_27 ( BL27, BLN27, WL15);
sram_cell_6t_3 inst_cell_15_26 ( BL26, BLN26, WL15);
sram_cell_6t_3 inst_cell_15_25 ( BL25, BLN25, WL15);
sram_cell_6t_3 inst_cell_15_24 ( BL24, BLN24, WL15);
sram_cell_6t_3 inst_cell_15_23 ( BL23, BLN23, WL15);
sram_cell_6t_3 inst_cell_15_22 ( BL22, BLN22, WL15);
sram_cell_6t_3 inst_cell_15_21 ( BL21, BLN21, WL15);
sram_cell_6t_3 inst_cell_15_20 ( BL20, BLN20, WL15);
sram_cell_6t_3 inst_cell_15_19 ( BL19, BLN19, WL15);
sram_cell_6t_3 inst_cell_15_18 ( BL18, BLN18, WL15);
sram_cell_6t_3 inst_cell_15_17 ( BL17, BLN17, WL15);
sram_cell_6t_3 inst_cell_15_16 ( BL16, BLN16, WL15);
sram_cell_6t_3 inst_cell_15_15 ( BL15, BLN15, WL15);
sram_cell_6t_3 inst_cell_15_14 ( BL14, BLN14, WL15);
sram_cell_6t_3 inst_cell_15_13 ( BL13, BLN13, WL15);
sram_cell_6t_3 inst_cell_15_12 ( BL12, BLN12, WL15);
sram_cell_6t_3 inst_cell_15_11 ( BL11, BLN11, WL15);
sram_cell_6t_3 inst_cell_15_10 ( BL10, BLN10, WL15);
sram_cell_6t_3 inst_cell_15_9 ( BL9, BLN9, WL15);
sram_cell_6t_3 inst_cell_15_8 ( BL8, BLN8, WL15);
sram_cell_6t_3 inst_cell_15_7 ( BL7, BLN7, WL15);
sram_cell_6t_3 inst_cell_15_6 ( BL6, BLN6, WL15);
sram_cell_6t_3 inst_cell_15_5 ( BL5, BLN5, WL15);
sram_cell_6t_3 inst_cell_15_4 ( BL4, BLN4, WL15);
sram_cell_6t_3 inst_cell_15_3 ( BL3, BLN3, WL15);
sram_cell_6t_3 inst_cell_15_2 ( BL2, BLN2, WL15);
sram_cell_6t_3 inst_cell_15_1 ( BL1, BLN1, WL15);
sram_cell_6t_3 inst_cell_15_0 ( BL0, BLN0, WL15);
sram_cell_6t_3 inst_cell_14_127 ( BL127, BLN127, WL14);
sram_cell_6t_3 inst_cell_14_126 ( BL126, BLN126, WL14);
sram_cell_6t_3 inst_cell_14_125 ( BL125, BLN125, WL14);
sram_cell_6t_3 inst_cell_14_124 ( BL124, BLN124, WL14);
sram_cell_6t_3 inst_cell_14_123 ( BL123, BLN123, WL14);
sram_cell_6t_3 inst_cell_14_122 ( BL122, BLN122, WL14);
sram_cell_6t_3 inst_cell_14_121 ( BL121, BLN121, WL14);
sram_cell_6t_3 inst_cell_14_120 ( BL120, BLN120, WL14);
sram_cell_6t_3 inst_cell_14_119 ( BL119, BLN119, WL14);
sram_cell_6t_3 inst_cell_14_118 ( BL118, BLN118, WL14);
sram_cell_6t_3 inst_cell_14_117 ( BL117, BLN117, WL14);
sram_cell_6t_3 inst_cell_14_116 ( BL116, BLN116, WL14);
sram_cell_6t_3 inst_cell_14_115 ( BL115, BLN115, WL14);
sram_cell_6t_3 inst_cell_14_114 ( BL114, BLN114, WL14);
sram_cell_6t_3 inst_cell_14_113 ( BL113, BLN113, WL14);
sram_cell_6t_3 inst_cell_14_112 ( BL112, BLN112, WL14);
sram_cell_6t_3 inst_cell_14_111 ( BL111, BLN111, WL14);
sram_cell_6t_3 inst_cell_14_110 ( BL110, BLN110, WL14);
sram_cell_6t_3 inst_cell_14_109 ( BL109, BLN109, WL14);
sram_cell_6t_3 inst_cell_14_108 ( BL108, BLN108, WL14);
sram_cell_6t_3 inst_cell_14_107 ( BL107, BLN107, WL14);
sram_cell_6t_3 inst_cell_14_106 ( BL106, BLN106, WL14);
sram_cell_6t_3 inst_cell_14_105 ( BL105, BLN105, WL14);
sram_cell_6t_3 inst_cell_14_104 ( BL104, BLN104, WL14);
sram_cell_6t_3 inst_cell_14_103 ( BL103, BLN103, WL14);
sram_cell_6t_3 inst_cell_14_102 ( BL102, BLN102, WL14);
sram_cell_6t_3 inst_cell_14_101 ( BL101, BLN101, WL14);
sram_cell_6t_3 inst_cell_14_100 ( BL100, BLN100, WL14);
sram_cell_6t_3 inst_cell_14_99 ( BL99, BLN99, WL14);
sram_cell_6t_3 inst_cell_14_98 ( BL98, BLN98, WL14);
sram_cell_6t_3 inst_cell_14_97 ( BL97, BLN97, WL14);
sram_cell_6t_3 inst_cell_14_96 ( BL96, BLN96, WL14);
sram_cell_6t_3 inst_cell_14_95 ( BL95, BLN95, WL14);
sram_cell_6t_3 inst_cell_14_94 ( BL94, BLN94, WL14);
sram_cell_6t_3 inst_cell_14_93 ( BL93, BLN93, WL14);
sram_cell_6t_3 inst_cell_14_92 ( BL92, BLN92, WL14);
sram_cell_6t_3 inst_cell_14_91 ( BL91, BLN91, WL14);
sram_cell_6t_3 inst_cell_14_90 ( BL90, BLN90, WL14);
sram_cell_6t_3 inst_cell_14_89 ( BL89, BLN89, WL14);
sram_cell_6t_3 inst_cell_14_88 ( BL88, BLN88, WL14);
sram_cell_6t_3 inst_cell_14_87 ( BL87, BLN87, WL14);
sram_cell_6t_3 inst_cell_14_86 ( BL86, BLN86, WL14);
sram_cell_6t_3 inst_cell_14_85 ( BL85, BLN85, WL14);
sram_cell_6t_3 inst_cell_14_84 ( BL84, BLN84, WL14);
sram_cell_6t_3 inst_cell_14_83 ( BL83, BLN83, WL14);
sram_cell_6t_3 inst_cell_14_82 ( BL82, BLN82, WL14);
sram_cell_6t_3 inst_cell_14_81 ( BL81, BLN81, WL14);
sram_cell_6t_3 inst_cell_14_80 ( BL80, BLN80, WL14);
sram_cell_6t_3 inst_cell_14_79 ( BL79, BLN79, WL14);
sram_cell_6t_3 inst_cell_14_78 ( BL78, BLN78, WL14);
sram_cell_6t_3 inst_cell_14_77 ( BL77, BLN77, WL14);
sram_cell_6t_3 inst_cell_14_76 ( BL76, BLN76, WL14);
sram_cell_6t_3 inst_cell_14_75 ( BL75, BLN75, WL14);
sram_cell_6t_3 inst_cell_14_74 ( BL74, BLN74, WL14);
sram_cell_6t_3 inst_cell_14_73 ( BL73, BLN73, WL14);
sram_cell_6t_3 inst_cell_14_72 ( BL72, BLN72, WL14);
sram_cell_6t_3 inst_cell_14_71 ( BL71, BLN71, WL14);
sram_cell_6t_3 inst_cell_14_70 ( BL70, BLN70, WL14);
sram_cell_6t_3 inst_cell_14_69 ( BL69, BLN69, WL14);
sram_cell_6t_3 inst_cell_14_68 ( BL68, BLN68, WL14);
sram_cell_6t_3 inst_cell_14_67 ( BL67, BLN67, WL14);
sram_cell_6t_3 inst_cell_14_66 ( BL66, BLN66, WL14);
sram_cell_6t_3 inst_cell_14_65 ( BL65, BLN65, WL14);
sram_cell_6t_3 inst_cell_14_64 ( BL64, BLN64, WL14);
sram_cell_6t_3 inst_cell_14_63 ( BL63, BLN63, WL14);
sram_cell_6t_3 inst_cell_14_62 ( BL62, BLN62, WL14);
sram_cell_6t_3 inst_cell_14_61 ( BL61, BLN61, WL14);
sram_cell_6t_3 inst_cell_14_60 ( BL60, BLN60, WL14);
sram_cell_6t_3 inst_cell_14_59 ( BL59, BLN59, WL14);
sram_cell_6t_3 inst_cell_14_58 ( BL58, BLN58, WL14);
sram_cell_6t_3 inst_cell_14_57 ( BL57, BLN57, WL14);
sram_cell_6t_3 inst_cell_14_56 ( BL56, BLN56, WL14);
sram_cell_6t_3 inst_cell_14_55 ( BL55, BLN55, WL14);
sram_cell_6t_3 inst_cell_14_54 ( BL54, BLN54, WL14);
sram_cell_6t_3 inst_cell_14_53 ( BL53, BLN53, WL14);
sram_cell_6t_3 inst_cell_14_52 ( BL52, BLN52, WL14);
sram_cell_6t_3 inst_cell_14_51 ( BL51, BLN51, WL14);
sram_cell_6t_3 inst_cell_14_50 ( BL50, BLN50, WL14);
sram_cell_6t_3 inst_cell_14_49 ( BL49, BLN49, WL14);
sram_cell_6t_3 inst_cell_14_48 ( BL48, BLN48, WL14);
sram_cell_6t_3 inst_cell_14_47 ( BL47, BLN47, WL14);
sram_cell_6t_3 inst_cell_14_46 ( BL46, BLN46, WL14);
sram_cell_6t_3 inst_cell_14_45 ( BL45, BLN45, WL14);
sram_cell_6t_3 inst_cell_14_44 ( BL44, BLN44, WL14);
sram_cell_6t_3 inst_cell_14_43 ( BL43, BLN43, WL14);
sram_cell_6t_3 inst_cell_14_42 ( BL42, BLN42, WL14);
sram_cell_6t_3 inst_cell_14_41 ( BL41, BLN41, WL14);
sram_cell_6t_3 inst_cell_14_40 ( BL40, BLN40, WL14);
sram_cell_6t_3 inst_cell_14_39 ( BL39, BLN39, WL14);
sram_cell_6t_3 inst_cell_14_38 ( BL38, BLN38, WL14);
sram_cell_6t_3 inst_cell_14_37 ( BL37, BLN37, WL14);
sram_cell_6t_3 inst_cell_14_36 ( BL36, BLN36, WL14);
sram_cell_6t_3 inst_cell_14_35 ( BL35, BLN35, WL14);
sram_cell_6t_3 inst_cell_14_34 ( BL34, BLN34, WL14);
sram_cell_6t_3 inst_cell_14_33 ( BL33, BLN33, WL14);
sram_cell_6t_3 inst_cell_14_32 ( BL32, BLN32, WL14);
sram_cell_6t_3 inst_cell_14_31 ( BL31, BLN31, WL14);
sram_cell_6t_3 inst_cell_14_30 ( BL30, BLN30, WL14);
sram_cell_6t_3 inst_cell_14_29 ( BL29, BLN29, WL14);
sram_cell_6t_3 inst_cell_14_28 ( BL28, BLN28, WL14);
sram_cell_6t_3 inst_cell_14_27 ( BL27, BLN27, WL14);
sram_cell_6t_3 inst_cell_14_26 ( BL26, BLN26, WL14);
sram_cell_6t_3 inst_cell_14_25 ( BL25, BLN25, WL14);
sram_cell_6t_3 inst_cell_14_24 ( BL24, BLN24, WL14);
sram_cell_6t_3 inst_cell_14_23 ( BL23, BLN23, WL14);
sram_cell_6t_3 inst_cell_14_22 ( BL22, BLN22, WL14);
sram_cell_6t_3 inst_cell_14_21 ( BL21, BLN21, WL14);
sram_cell_6t_3 inst_cell_14_20 ( BL20, BLN20, WL14);
sram_cell_6t_3 inst_cell_14_19 ( BL19, BLN19, WL14);
sram_cell_6t_3 inst_cell_14_18 ( BL18, BLN18, WL14);
sram_cell_6t_3 inst_cell_14_17 ( BL17, BLN17, WL14);
sram_cell_6t_3 inst_cell_14_16 ( BL16, BLN16, WL14);
sram_cell_6t_3 inst_cell_14_15 ( BL15, BLN15, WL14);
sram_cell_6t_3 inst_cell_14_14 ( BL14, BLN14, WL14);
sram_cell_6t_3 inst_cell_14_13 ( BL13, BLN13, WL14);
sram_cell_6t_3 inst_cell_14_12 ( BL12, BLN12, WL14);
sram_cell_6t_3 inst_cell_14_11 ( BL11, BLN11, WL14);
sram_cell_6t_3 inst_cell_14_10 ( BL10, BLN10, WL14);
sram_cell_6t_3 inst_cell_14_9 ( BL9, BLN9, WL14);
sram_cell_6t_3 inst_cell_14_8 ( BL8, BLN8, WL14);
sram_cell_6t_3 inst_cell_14_7 ( BL7, BLN7, WL14);
sram_cell_6t_3 inst_cell_14_6 ( BL6, BLN6, WL14);
sram_cell_6t_3 inst_cell_14_5 ( BL5, BLN5, WL14);
sram_cell_6t_3 inst_cell_14_4 ( BL4, BLN4, WL14);
sram_cell_6t_3 inst_cell_14_3 ( BL3, BLN3, WL14);
sram_cell_6t_3 inst_cell_14_2 ( BL2, BLN2, WL14);
sram_cell_6t_3 inst_cell_14_1 ( BL1, BLN1, WL14);
sram_cell_6t_3 inst_cell_14_0 ( BL0, BLN0, WL14);
sram_cell_6t_3 inst_cell_13_127 ( BL127, BLN127, WL13);
sram_cell_6t_3 inst_cell_12_127 ( BL127, BLN127, WL12);
sram_cell_6t_3 inst_cell_11_127 ( BL127, BLN127, WL11);
sram_cell_6t_3 inst_cell_10_127 ( BL127, BLN127, WL10);
sram_cell_6t_3 inst_cell_9_127 ( BL127, BLN127, WL9);
sram_cell_6t_3 inst_cell_8_127 ( BL127, BLN127, WL8);
sram_cell_6t_3 inst_cell_7_127 ( BL127, BLN127, WL7);
sram_cell_6t_3 inst_cell_6_127 ( BL127, BLN127, WL6);
sram_cell_6t_3 inst_cell_5_127 ( BL127, BLN127, WL5);
sram_cell_6t_3 inst_cell_4_127 ( BL127, BLN127, WL4);
sram_cell_6t_3 inst_cell_3_127 ( BL127, BLN127, WL3);
sram_cell_6t_3 inst_cell_2_127 ( BL127, BLN127, WL2);
sram_cell_6t_3 inst_cell_1_127 ( BL127, BLN127, WL1);
sram_cell_6t_3 inst_cell_0_127 ( BL127, BLN127, WL0);
sram_cell_6t_3 inst_cell_13_126 ( BL126, BLN126, WL13);
sram_cell_6t_3 inst_cell_12_126 ( BL126, BLN126, WL12);
sram_cell_6t_3 inst_cell_11_126 ( BL126, BLN126, WL11);
sram_cell_6t_3 inst_cell_10_126 ( BL126, BLN126, WL10);
sram_cell_6t_3 inst_cell_9_126 ( BL126, BLN126, WL9);
sram_cell_6t_3 inst_cell_8_126 ( BL126, BLN126, WL8);
sram_cell_6t_3 inst_cell_7_126 ( BL126, BLN126, WL7);
sram_cell_6t_3 inst_cell_6_126 ( BL126, BLN126, WL6);
sram_cell_6t_3 inst_cell_5_126 ( BL126, BLN126, WL5);
sram_cell_6t_3 inst_cell_4_126 ( BL126, BLN126, WL4);
sram_cell_6t_3 inst_cell_3_126 ( BL126, BLN126, WL3);
sram_cell_6t_3 inst_cell_2_126 ( BL126, BLN126, WL2);
sram_cell_6t_3 inst_cell_1_126 ( BL126, BLN126, WL1);
sram_cell_6t_3 inst_cell_0_126 ( BL126, BLN126, WL0);
sram_cell_6t_3 inst_cell_13_125 ( BL125, BLN125, WL13);
sram_cell_6t_3 inst_cell_12_125 ( BL125, BLN125, WL12);
sram_cell_6t_3 inst_cell_11_125 ( BL125, BLN125, WL11);
sram_cell_6t_3 inst_cell_10_125 ( BL125, BLN125, WL10);
sram_cell_6t_3 inst_cell_9_125 ( BL125, BLN125, WL9);
sram_cell_6t_3 inst_cell_8_125 ( BL125, BLN125, WL8);
sram_cell_6t_3 inst_cell_7_125 ( BL125, BLN125, WL7);
sram_cell_6t_3 inst_cell_6_125 ( BL125, BLN125, WL6);
sram_cell_6t_3 inst_cell_5_125 ( BL125, BLN125, WL5);
sram_cell_6t_3 inst_cell_4_125 ( BL125, BLN125, WL4);
sram_cell_6t_3 inst_cell_3_125 ( BL125, BLN125, WL3);
sram_cell_6t_3 inst_cell_2_125 ( BL125, BLN125, WL2);
sram_cell_6t_3 inst_cell_1_125 ( BL125, BLN125, WL1);
sram_cell_6t_3 inst_cell_0_125 ( BL125, BLN125, WL0);
sram_cell_6t_3 inst_cell_13_124 ( BL124, BLN124, WL13);
sram_cell_6t_3 inst_cell_12_124 ( BL124, BLN124, WL12);
sram_cell_6t_3 inst_cell_11_124 ( BL124, BLN124, WL11);
sram_cell_6t_3 inst_cell_10_124 ( BL124, BLN124, WL10);
sram_cell_6t_3 inst_cell_9_124 ( BL124, BLN124, WL9);
sram_cell_6t_3 inst_cell_8_124 ( BL124, BLN124, WL8);
sram_cell_6t_3 inst_cell_7_124 ( BL124, BLN124, WL7);
sram_cell_6t_3 inst_cell_6_124 ( BL124, BLN124, WL6);
sram_cell_6t_3 inst_cell_5_124 ( BL124, BLN124, WL5);
sram_cell_6t_3 inst_cell_4_124 ( BL124, BLN124, WL4);
sram_cell_6t_3 inst_cell_3_124 ( BL124, BLN124, WL3);
sram_cell_6t_3 inst_cell_2_124 ( BL124, BLN124, WL2);
sram_cell_6t_3 inst_cell_1_124 ( BL124, BLN124, WL1);
sram_cell_6t_3 inst_cell_0_124 ( BL124, BLN124, WL0);
sram_cell_6t_3 inst_cell_13_123 ( BL123, BLN123, WL13);
sram_cell_6t_3 inst_cell_12_123 ( BL123, BLN123, WL12);
sram_cell_6t_3 inst_cell_11_123 ( BL123, BLN123, WL11);
sram_cell_6t_3 inst_cell_10_123 ( BL123, BLN123, WL10);
sram_cell_6t_3 inst_cell_9_123 ( BL123, BLN123, WL9);
sram_cell_6t_3 inst_cell_8_123 ( BL123, BLN123, WL8);
sram_cell_6t_3 inst_cell_7_123 ( BL123, BLN123, WL7);
sram_cell_6t_3 inst_cell_6_123 ( BL123, BLN123, WL6);
sram_cell_6t_3 inst_cell_5_123 ( BL123, BLN123, WL5);
sram_cell_6t_3 inst_cell_4_123 ( BL123, BLN123, WL4);
sram_cell_6t_3 inst_cell_3_123 ( BL123, BLN123, WL3);
sram_cell_6t_3 inst_cell_2_123 ( BL123, BLN123, WL2);
sram_cell_6t_3 inst_cell_1_123 ( BL123, BLN123, WL1);
sram_cell_6t_3 inst_cell_0_123 ( BL123, BLN123, WL0);
sram_cell_6t_3 inst_cell_13_122 ( BL122, BLN122, WL13);
sram_cell_6t_3 inst_cell_12_122 ( BL122, BLN122, WL12);
sram_cell_6t_3 inst_cell_11_122 ( BL122, BLN122, WL11);
sram_cell_6t_3 inst_cell_10_122 ( BL122, BLN122, WL10);
sram_cell_6t_3 inst_cell_9_122 ( BL122, BLN122, WL9);
sram_cell_6t_3 inst_cell_8_122 ( BL122, BLN122, WL8);
sram_cell_6t_3 inst_cell_7_122 ( BL122, BLN122, WL7);
sram_cell_6t_3 inst_cell_6_122 ( BL122, BLN122, WL6);
sram_cell_6t_3 inst_cell_5_122 ( BL122, BLN122, WL5);
sram_cell_6t_3 inst_cell_4_122 ( BL122, BLN122, WL4);
sram_cell_6t_3 inst_cell_3_122 ( BL122, BLN122, WL3);
sram_cell_6t_3 inst_cell_2_122 ( BL122, BLN122, WL2);
sram_cell_6t_3 inst_cell_1_122 ( BL122, BLN122, WL1);
sram_cell_6t_3 inst_cell_0_122 ( BL122, BLN122, WL0);
sram_cell_6t_3 inst_cell_13_121 ( BL121, BLN121, WL13);
sram_cell_6t_3 inst_cell_12_121 ( BL121, BLN121, WL12);
sram_cell_6t_3 inst_cell_11_121 ( BL121, BLN121, WL11);
sram_cell_6t_3 inst_cell_10_121 ( BL121, BLN121, WL10);
sram_cell_6t_3 inst_cell_9_121 ( BL121, BLN121, WL9);
sram_cell_6t_3 inst_cell_8_121 ( BL121, BLN121, WL8);
sram_cell_6t_3 inst_cell_7_121 ( BL121, BLN121, WL7);
sram_cell_6t_3 inst_cell_6_121 ( BL121, BLN121, WL6);
sram_cell_6t_3 inst_cell_5_121 ( BL121, BLN121, WL5);
sram_cell_6t_3 inst_cell_4_121 ( BL121, BLN121, WL4);
sram_cell_6t_3 inst_cell_3_121 ( BL121, BLN121, WL3);
sram_cell_6t_3 inst_cell_2_121 ( BL121, BLN121, WL2);
sram_cell_6t_3 inst_cell_1_121 ( BL121, BLN121, WL1);
sram_cell_6t_3 inst_cell_0_121 ( BL121, BLN121, WL0);
sram_cell_6t_3 inst_cell_13_120 ( BL120, BLN120, WL13);
sram_cell_6t_3 inst_cell_12_120 ( BL120, BLN120, WL12);
sram_cell_6t_3 inst_cell_11_120 ( BL120, BLN120, WL11);
sram_cell_6t_3 inst_cell_10_120 ( BL120, BLN120, WL10);
sram_cell_6t_3 inst_cell_9_120 ( BL120, BLN120, WL9);
sram_cell_6t_3 inst_cell_8_120 ( BL120, BLN120, WL8);
sram_cell_6t_3 inst_cell_7_120 ( BL120, BLN120, WL7);
sram_cell_6t_3 inst_cell_6_120 ( BL120, BLN120, WL6);
sram_cell_6t_3 inst_cell_5_120 ( BL120, BLN120, WL5);
sram_cell_6t_3 inst_cell_4_120 ( BL120, BLN120, WL4);
sram_cell_6t_3 inst_cell_3_120 ( BL120, BLN120, WL3);
sram_cell_6t_3 inst_cell_2_120 ( BL120, BLN120, WL2);
sram_cell_6t_3 inst_cell_1_120 ( BL120, BLN120, WL1);
sram_cell_6t_3 inst_cell_0_120 ( BL120, BLN120, WL0);
sram_cell_6t_3 inst_cell_13_119 ( BL119, BLN119, WL13);
sram_cell_6t_3 inst_cell_12_119 ( BL119, BLN119, WL12);
sram_cell_6t_3 inst_cell_11_119 ( BL119, BLN119, WL11);
sram_cell_6t_3 inst_cell_10_119 ( BL119, BLN119, WL10);
sram_cell_6t_3 inst_cell_9_119 ( BL119, BLN119, WL9);
sram_cell_6t_3 inst_cell_8_119 ( BL119, BLN119, WL8);
sram_cell_6t_3 inst_cell_7_119 ( BL119, BLN119, WL7);
sram_cell_6t_3 inst_cell_6_119 ( BL119, BLN119, WL6);
sram_cell_6t_3 inst_cell_5_119 ( BL119, BLN119, WL5);
sram_cell_6t_3 inst_cell_4_119 ( BL119, BLN119, WL4);
sram_cell_6t_3 inst_cell_3_119 ( BL119, BLN119, WL3);
sram_cell_6t_3 inst_cell_2_119 ( BL119, BLN119, WL2);
sram_cell_6t_3 inst_cell_1_119 ( BL119, BLN119, WL1);
sram_cell_6t_3 inst_cell_0_119 ( BL119, BLN119, WL0);
sram_cell_6t_3 inst_cell_13_118 ( BL118, BLN118, WL13);
sram_cell_6t_3 inst_cell_12_118 ( BL118, BLN118, WL12);
sram_cell_6t_3 inst_cell_11_118 ( BL118, BLN118, WL11);
sram_cell_6t_3 inst_cell_10_118 ( BL118, BLN118, WL10);
sram_cell_6t_3 inst_cell_9_118 ( BL118, BLN118, WL9);
sram_cell_6t_3 inst_cell_8_118 ( BL118, BLN118, WL8);
sram_cell_6t_3 inst_cell_7_118 ( BL118, BLN118, WL7);
sram_cell_6t_3 inst_cell_6_118 ( BL118, BLN118, WL6);
sram_cell_6t_3 inst_cell_5_118 ( BL118, BLN118, WL5);
sram_cell_6t_3 inst_cell_4_118 ( BL118, BLN118, WL4);
sram_cell_6t_3 inst_cell_3_118 ( BL118, BLN118, WL3);
sram_cell_6t_3 inst_cell_2_118 ( BL118, BLN118, WL2);
sram_cell_6t_3 inst_cell_1_118 ( BL118, BLN118, WL1);
sram_cell_6t_3 inst_cell_0_118 ( BL118, BLN118, WL0);
sram_cell_6t_3 inst_cell_13_117 ( BL117, BLN117, WL13);
sram_cell_6t_3 inst_cell_12_117 ( BL117, BLN117, WL12);
sram_cell_6t_3 inst_cell_11_117 ( BL117, BLN117, WL11);
sram_cell_6t_3 inst_cell_10_117 ( BL117, BLN117, WL10);
sram_cell_6t_3 inst_cell_9_117 ( BL117, BLN117, WL9);
sram_cell_6t_3 inst_cell_8_117 ( BL117, BLN117, WL8);
sram_cell_6t_3 inst_cell_7_117 ( BL117, BLN117, WL7);
sram_cell_6t_3 inst_cell_6_117 ( BL117, BLN117, WL6);
sram_cell_6t_3 inst_cell_5_117 ( BL117, BLN117, WL5);
sram_cell_6t_3 inst_cell_4_117 ( BL117, BLN117, WL4);
sram_cell_6t_3 inst_cell_3_117 ( BL117, BLN117, WL3);
sram_cell_6t_3 inst_cell_2_117 ( BL117, BLN117, WL2);
sram_cell_6t_3 inst_cell_1_117 ( BL117, BLN117, WL1);
sram_cell_6t_3 inst_cell_0_117 ( BL117, BLN117, WL0);
sram_cell_6t_3 inst_cell_13_116 ( BL116, BLN116, WL13);
sram_cell_6t_3 inst_cell_12_116 ( BL116, BLN116, WL12);
sram_cell_6t_3 inst_cell_11_116 ( BL116, BLN116, WL11);
sram_cell_6t_3 inst_cell_10_116 ( BL116, BLN116, WL10);
sram_cell_6t_3 inst_cell_9_116 ( BL116, BLN116, WL9);
sram_cell_6t_3 inst_cell_8_116 ( BL116, BLN116, WL8);
sram_cell_6t_3 inst_cell_7_116 ( BL116, BLN116, WL7);
sram_cell_6t_3 inst_cell_6_116 ( BL116, BLN116, WL6);
sram_cell_6t_3 inst_cell_5_116 ( BL116, BLN116, WL5);
sram_cell_6t_3 inst_cell_4_116 ( BL116, BLN116, WL4);
sram_cell_6t_3 inst_cell_3_116 ( BL116, BLN116, WL3);
sram_cell_6t_3 inst_cell_2_116 ( BL116, BLN116, WL2);
sram_cell_6t_3 inst_cell_1_116 ( BL116, BLN116, WL1);
sram_cell_6t_3 inst_cell_0_116 ( BL116, BLN116, WL0);
sram_cell_6t_3 inst_cell_13_115 ( BL115, BLN115, WL13);
sram_cell_6t_3 inst_cell_12_115 ( BL115, BLN115, WL12);
sram_cell_6t_3 inst_cell_11_115 ( BL115, BLN115, WL11);
sram_cell_6t_3 inst_cell_10_115 ( BL115, BLN115, WL10);
sram_cell_6t_3 inst_cell_9_115 ( BL115, BLN115, WL9);
sram_cell_6t_3 inst_cell_8_115 ( BL115, BLN115, WL8);
sram_cell_6t_3 inst_cell_7_115 ( BL115, BLN115, WL7);
sram_cell_6t_3 inst_cell_6_115 ( BL115, BLN115, WL6);
sram_cell_6t_3 inst_cell_5_115 ( BL115, BLN115, WL5);
sram_cell_6t_3 inst_cell_4_115 ( BL115, BLN115, WL4);
sram_cell_6t_3 inst_cell_3_115 ( BL115, BLN115, WL3);
sram_cell_6t_3 inst_cell_2_115 ( BL115, BLN115, WL2);
sram_cell_6t_3 inst_cell_1_115 ( BL115, BLN115, WL1);
sram_cell_6t_3 inst_cell_0_115 ( BL115, BLN115, WL0);
sram_cell_6t_3 inst_cell_13_114 ( BL114, BLN114, WL13);
sram_cell_6t_3 inst_cell_12_114 ( BL114, BLN114, WL12);
sram_cell_6t_3 inst_cell_11_114 ( BL114, BLN114, WL11);
sram_cell_6t_3 inst_cell_10_114 ( BL114, BLN114, WL10);
sram_cell_6t_3 inst_cell_9_114 ( BL114, BLN114, WL9);
sram_cell_6t_3 inst_cell_8_114 ( BL114, BLN114, WL8);
sram_cell_6t_3 inst_cell_7_114 ( BL114, BLN114, WL7);
sram_cell_6t_3 inst_cell_6_114 ( BL114, BLN114, WL6);
sram_cell_6t_3 inst_cell_5_114 ( BL114, BLN114, WL5);
sram_cell_6t_3 inst_cell_4_114 ( BL114, BLN114, WL4);
sram_cell_6t_3 inst_cell_3_114 ( BL114, BLN114, WL3);
sram_cell_6t_3 inst_cell_2_114 ( BL114, BLN114, WL2);
sram_cell_6t_3 inst_cell_1_114 ( BL114, BLN114, WL1);
sram_cell_6t_3 inst_cell_0_114 ( BL114, BLN114, WL0);
sram_cell_6t_3 inst_cell_13_113 ( BL113, BLN113, WL13);
sram_cell_6t_3 inst_cell_12_113 ( BL113, BLN113, WL12);
sram_cell_6t_3 inst_cell_11_113 ( BL113, BLN113, WL11);
sram_cell_6t_3 inst_cell_10_113 ( BL113, BLN113, WL10);
sram_cell_6t_3 inst_cell_9_113 ( BL113, BLN113, WL9);
sram_cell_6t_3 inst_cell_8_113 ( BL113, BLN113, WL8);
sram_cell_6t_3 inst_cell_7_113 ( BL113, BLN113, WL7);
sram_cell_6t_3 inst_cell_6_113 ( BL113, BLN113, WL6);
sram_cell_6t_3 inst_cell_5_113 ( BL113, BLN113, WL5);
sram_cell_6t_3 inst_cell_4_113 ( BL113, BLN113, WL4);
sram_cell_6t_3 inst_cell_3_113 ( BL113, BLN113, WL3);
sram_cell_6t_3 inst_cell_2_113 ( BL113, BLN113, WL2);
sram_cell_6t_3 inst_cell_1_113 ( BL113, BLN113, WL1);
sram_cell_6t_3 inst_cell_0_113 ( BL113, BLN113, WL0);
sram_cell_6t_3 inst_cell_13_112 ( BL112, BLN112, WL13);
sram_cell_6t_3 inst_cell_12_112 ( BL112, BLN112, WL12);
sram_cell_6t_3 inst_cell_11_112 ( BL112, BLN112, WL11);
sram_cell_6t_3 inst_cell_10_112 ( BL112, BLN112, WL10);
sram_cell_6t_3 inst_cell_9_112 ( BL112, BLN112, WL9);
sram_cell_6t_3 inst_cell_8_112 ( BL112, BLN112, WL8);
sram_cell_6t_3 inst_cell_7_112 ( BL112, BLN112, WL7);
sram_cell_6t_3 inst_cell_6_112 ( BL112, BLN112, WL6);
sram_cell_6t_3 inst_cell_5_112 ( BL112, BLN112, WL5);
sram_cell_6t_3 inst_cell_4_112 ( BL112, BLN112, WL4);
sram_cell_6t_3 inst_cell_3_112 ( BL112, BLN112, WL3);
sram_cell_6t_3 inst_cell_2_112 ( BL112, BLN112, WL2);
sram_cell_6t_3 inst_cell_1_112 ( BL112, BLN112, WL1);
sram_cell_6t_3 inst_cell_0_112 ( BL112, BLN112, WL0);
sram_cell_6t_3 inst_cell_13_111 ( BL111, BLN111, WL13);
sram_cell_6t_3 inst_cell_12_111 ( BL111, BLN111, WL12);
sram_cell_6t_3 inst_cell_11_111 ( BL111, BLN111, WL11);
sram_cell_6t_3 inst_cell_10_111 ( BL111, BLN111, WL10);
sram_cell_6t_3 inst_cell_9_111 ( BL111, BLN111, WL9);
sram_cell_6t_3 inst_cell_8_111 ( BL111, BLN111, WL8);
sram_cell_6t_3 inst_cell_7_111 ( BL111, BLN111, WL7);
sram_cell_6t_3 inst_cell_6_111 ( BL111, BLN111, WL6);
sram_cell_6t_3 inst_cell_5_111 ( BL111, BLN111, WL5);
sram_cell_6t_3 inst_cell_4_111 ( BL111, BLN111, WL4);
sram_cell_6t_3 inst_cell_3_111 ( BL111, BLN111, WL3);
sram_cell_6t_3 inst_cell_2_111 ( BL111, BLN111, WL2);
sram_cell_6t_3 inst_cell_1_111 ( BL111, BLN111, WL1);
sram_cell_6t_3 inst_cell_0_111 ( BL111, BLN111, WL0);
sram_cell_6t_3 inst_cell_13_110 ( BL110, BLN110, WL13);
sram_cell_6t_3 inst_cell_12_110 ( BL110, BLN110, WL12);
sram_cell_6t_3 inst_cell_11_110 ( BL110, BLN110, WL11);
sram_cell_6t_3 inst_cell_10_110 ( BL110, BLN110, WL10);
sram_cell_6t_3 inst_cell_9_110 ( BL110, BLN110, WL9);
sram_cell_6t_3 inst_cell_8_110 ( BL110, BLN110, WL8);
sram_cell_6t_3 inst_cell_7_110 ( BL110, BLN110, WL7);
sram_cell_6t_3 inst_cell_6_110 ( BL110, BLN110, WL6);
sram_cell_6t_3 inst_cell_5_110 ( BL110, BLN110, WL5);
sram_cell_6t_3 inst_cell_4_110 ( BL110, BLN110, WL4);
sram_cell_6t_3 inst_cell_3_110 ( BL110, BLN110, WL3);
sram_cell_6t_3 inst_cell_2_110 ( BL110, BLN110, WL2);
sram_cell_6t_3 inst_cell_1_110 ( BL110, BLN110, WL1);
sram_cell_6t_3 inst_cell_0_110 ( BL110, BLN110, WL0);
sram_cell_6t_3 inst_cell_13_109 ( BL109, BLN109, WL13);
sram_cell_6t_3 inst_cell_12_109 ( BL109, BLN109, WL12);
sram_cell_6t_3 inst_cell_11_109 ( BL109, BLN109, WL11);
sram_cell_6t_3 inst_cell_10_109 ( BL109, BLN109, WL10);
sram_cell_6t_3 inst_cell_9_109 ( BL109, BLN109, WL9);
sram_cell_6t_3 inst_cell_8_109 ( BL109, BLN109, WL8);
sram_cell_6t_3 inst_cell_7_109 ( BL109, BLN109, WL7);
sram_cell_6t_3 inst_cell_6_109 ( BL109, BLN109, WL6);
sram_cell_6t_3 inst_cell_5_109 ( BL109, BLN109, WL5);
sram_cell_6t_3 inst_cell_4_109 ( BL109, BLN109, WL4);
sram_cell_6t_3 inst_cell_3_109 ( BL109, BLN109, WL3);
sram_cell_6t_3 inst_cell_2_109 ( BL109, BLN109, WL2);
sram_cell_6t_3 inst_cell_1_109 ( BL109, BLN109, WL1);
sram_cell_6t_3 inst_cell_0_109 ( BL109, BLN109, WL0);
sram_cell_6t_3 inst_cell_13_108 ( BL108, BLN108, WL13);
sram_cell_6t_3 inst_cell_12_108 ( BL108, BLN108, WL12);
sram_cell_6t_3 inst_cell_11_108 ( BL108, BLN108, WL11);
sram_cell_6t_3 inst_cell_10_108 ( BL108, BLN108, WL10);
sram_cell_6t_3 inst_cell_9_108 ( BL108, BLN108, WL9);
sram_cell_6t_3 inst_cell_8_108 ( BL108, BLN108, WL8);
sram_cell_6t_3 inst_cell_7_108 ( BL108, BLN108, WL7);
sram_cell_6t_3 inst_cell_6_108 ( BL108, BLN108, WL6);
sram_cell_6t_3 inst_cell_5_108 ( BL108, BLN108, WL5);
sram_cell_6t_3 inst_cell_4_108 ( BL108, BLN108, WL4);
sram_cell_6t_3 inst_cell_3_108 ( BL108, BLN108, WL3);
sram_cell_6t_3 inst_cell_2_108 ( BL108, BLN108, WL2);
sram_cell_6t_3 inst_cell_1_108 ( BL108, BLN108, WL1);
sram_cell_6t_3 inst_cell_0_108 ( BL108, BLN108, WL0);
sram_cell_6t_3 inst_cell_13_107 ( BL107, BLN107, WL13);
sram_cell_6t_3 inst_cell_12_107 ( BL107, BLN107, WL12);
sram_cell_6t_3 inst_cell_11_107 ( BL107, BLN107, WL11);
sram_cell_6t_3 inst_cell_10_107 ( BL107, BLN107, WL10);
sram_cell_6t_3 inst_cell_9_107 ( BL107, BLN107, WL9);
sram_cell_6t_3 inst_cell_8_107 ( BL107, BLN107, WL8);
sram_cell_6t_3 inst_cell_7_107 ( BL107, BLN107, WL7);
sram_cell_6t_3 inst_cell_6_107 ( BL107, BLN107, WL6);
sram_cell_6t_3 inst_cell_5_107 ( BL107, BLN107, WL5);
sram_cell_6t_3 inst_cell_4_107 ( BL107, BLN107, WL4);
sram_cell_6t_3 inst_cell_3_107 ( BL107, BLN107, WL3);
sram_cell_6t_3 inst_cell_2_107 ( BL107, BLN107, WL2);
sram_cell_6t_3 inst_cell_1_107 ( BL107, BLN107, WL1);
sram_cell_6t_3 inst_cell_0_107 ( BL107, BLN107, WL0);
sram_cell_6t_3 inst_cell_13_106 ( BL106, BLN106, WL13);
sram_cell_6t_3 inst_cell_12_106 ( BL106, BLN106, WL12);
sram_cell_6t_3 inst_cell_11_106 ( BL106, BLN106, WL11);
sram_cell_6t_3 inst_cell_10_106 ( BL106, BLN106, WL10);
sram_cell_6t_3 inst_cell_9_106 ( BL106, BLN106, WL9);
sram_cell_6t_3 inst_cell_8_106 ( BL106, BLN106, WL8);
sram_cell_6t_3 inst_cell_7_106 ( BL106, BLN106, WL7);
sram_cell_6t_3 inst_cell_6_106 ( BL106, BLN106, WL6);
sram_cell_6t_3 inst_cell_5_106 ( BL106, BLN106, WL5);
sram_cell_6t_3 inst_cell_4_106 ( BL106, BLN106, WL4);
sram_cell_6t_3 inst_cell_3_106 ( BL106, BLN106, WL3);
sram_cell_6t_3 inst_cell_2_106 ( BL106, BLN106, WL2);
sram_cell_6t_3 inst_cell_1_106 ( BL106, BLN106, WL1);
sram_cell_6t_3 inst_cell_0_106 ( BL106, BLN106, WL0);
sram_cell_6t_3 inst_cell_13_105 ( BL105, BLN105, WL13);
sram_cell_6t_3 inst_cell_12_105 ( BL105, BLN105, WL12);
sram_cell_6t_3 inst_cell_11_105 ( BL105, BLN105, WL11);
sram_cell_6t_3 inst_cell_10_105 ( BL105, BLN105, WL10);
sram_cell_6t_3 inst_cell_9_105 ( BL105, BLN105, WL9);
sram_cell_6t_3 inst_cell_8_105 ( BL105, BLN105, WL8);
sram_cell_6t_3 inst_cell_7_105 ( BL105, BLN105, WL7);
sram_cell_6t_3 inst_cell_6_105 ( BL105, BLN105, WL6);
sram_cell_6t_3 inst_cell_5_105 ( BL105, BLN105, WL5);
sram_cell_6t_3 inst_cell_4_105 ( BL105, BLN105, WL4);
sram_cell_6t_3 inst_cell_3_105 ( BL105, BLN105, WL3);
sram_cell_6t_3 inst_cell_2_105 ( BL105, BLN105, WL2);
sram_cell_6t_3 inst_cell_1_105 ( BL105, BLN105, WL1);
sram_cell_6t_3 inst_cell_0_105 ( BL105, BLN105, WL0);
sram_cell_6t_3 inst_cell_13_104 ( BL104, BLN104, WL13);
sram_cell_6t_3 inst_cell_12_104 ( BL104, BLN104, WL12);
sram_cell_6t_3 inst_cell_11_104 ( BL104, BLN104, WL11);
sram_cell_6t_3 inst_cell_10_104 ( BL104, BLN104, WL10);
sram_cell_6t_3 inst_cell_9_104 ( BL104, BLN104, WL9);
sram_cell_6t_3 inst_cell_8_104 ( BL104, BLN104, WL8);
sram_cell_6t_3 inst_cell_7_104 ( BL104, BLN104, WL7);
sram_cell_6t_3 inst_cell_6_104 ( BL104, BLN104, WL6);
sram_cell_6t_3 inst_cell_5_104 ( BL104, BLN104, WL5);
sram_cell_6t_3 inst_cell_4_104 ( BL104, BLN104, WL4);
sram_cell_6t_3 inst_cell_3_104 ( BL104, BLN104, WL3);
sram_cell_6t_3 inst_cell_2_104 ( BL104, BLN104, WL2);
sram_cell_6t_3 inst_cell_1_104 ( BL104, BLN104, WL1);
sram_cell_6t_3 inst_cell_0_104 ( BL104, BLN104, WL0);
sram_cell_6t_3 inst_cell_13_103 ( BL103, BLN103, WL13);
sram_cell_6t_3 inst_cell_12_103 ( BL103, BLN103, WL12);
sram_cell_6t_3 inst_cell_11_103 ( BL103, BLN103, WL11);
sram_cell_6t_3 inst_cell_10_103 ( BL103, BLN103, WL10);
sram_cell_6t_3 inst_cell_9_103 ( BL103, BLN103, WL9);
sram_cell_6t_3 inst_cell_8_103 ( BL103, BLN103, WL8);
sram_cell_6t_3 inst_cell_7_103 ( BL103, BLN103, WL7);
sram_cell_6t_3 inst_cell_6_103 ( BL103, BLN103, WL6);
sram_cell_6t_3 inst_cell_5_103 ( BL103, BLN103, WL5);
sram_cell_6t_3 inst_cell_4_103 ( BL103, BLN103, WL4);
sram_cell_6t_3 inst_cell_3_103 ( BL103, BLN103, WL3);
sram_cell_6t_3 inst_cell_2_103 ( BL103, BLN103, WL2);
sram_cell_6t_3 inst_cell_1_103 ( BL103, BLN103, WL1);
sram_cell_6t_3 inst_cell_0_103 ( BL103, BLN103, WL0);
sram_cell_6t_3 inst_cell_13_102 ( BL102, BLN102, WL13);
sram_cell_6t_3 inst_cell_12_102 ( BL102, BLN102, WL12);
sram_cell_6t_3 inst_cell_11_102 ( BL102, BLN102, WL11);
sram_cell_6t_3 inst_cell_10_102 ( BL102, BLN102, WL10);
sram_cell_6t_3 inst_cell_9_102 ( BL102, BLN102, WL9);
sram_cell_6t_3 inst_cell_8_102 ( BL102, BLN102, WL8);
sram_cell_6t_3 inst_cell_7_102 ( BL102, BLN102, WL7);
sram_cell_6t_3 inst_cell_6_102 ( BL102, BLN102, WL6);
sram_cell_6t_3 inst_cell_5_102 ( BL102, BLN102, WL5);
sram_cell_6t_3 inst_cell_4_102 ( BL102, BLN102, WL4);
sram_cell_6t_3 inst_cell_3_102 ( BL102, BLN102, WL3);
sram_cell_6t_3 inst_cell_2_102 ( BL102, BLN102, WL2);
sram_cell_6t_3 inst_cell_1_102 ( BL102, BLN102, WL1);
sram_cell_6t_3 inst_cell_0_102 ( BL102, BLN102, WL0);
sram_cell_6t_3 inst_cell_13_101 ( BL101, BLN101, WL13);
sram_cell_6t_3 inst_cell_12_101 ( BL101, BLN101, WL12);
sram_cell_6t_3 inst_cell_11_101 ( BL101, BLN101, WL11);
sram_cell_6t_3 inst_cell_10_101 ( BL101, BLN101, WL10);
sram_cell_6t_3 inst_cell_9_101 ( BL101, BLN101, WL9);
sram_cell_6t_3 inst_cell_8_101 ( BL101, BLN101, WL8);
sram_cell_6t_3 inst_cell_7_101 ( BL101, BLN101, WL7);
sram_cell_6t_3 inst_cell_6_101 ( BL101, BLN101, WL6);
sram_cell_6t_3 inst_cell_5_101 ( BL101, BLN101, WL5);
sram_cell_6t_3 inst_cell_4_101 ( BL101, BLN101, WL4);
sram_cell_6t_3 inst_cell_3_101 ( BL101, BLN101, WL3);
sram_cell_6t_3 inst_cell_2_101 ( BL101, BLN101, WL2);
sram_cell_6t_3 inst_cell_1_101 ( BL101, BLN101, WL1);
sram_cell_6t_3 inst_cell_0_101 ( BL101, BLN101, WL0);
sram_cell_6t_3 inst_cell_13_100 ( BL100, BLN100, WL13);
sram_cell_6t_3 inst_cell_12_100 ( BL100, BLN100, WL12);
sram_cell_6t_3 inst_cell_11_100 ( BL100, BLN100, WL11);
sram_cell_6t_3 inst_cell_10_100 ( BL100, BLN100, WL10);
sram_cell_6t_3 inst_cell_9_100 ( BL100, BLN100, WL9);
sram_cell_6t_3 inst_cell_8_100 ( BL100, BLN100, WL8);
sram_cell_6t_3 inst_cell_7_100 ( BL100, BLN100, WL7);
sram_cell_6t_3 inst_cell_6_100 ( BL100, BLN100, WL6);
sram_cell_6t_3 inst_cell_5_100 ( BL100, BLN100, WL5);
sram_cell_6t_3 inst_cell_4_100 ( BL100, BLN100, WL4);
sram_cell_6t_3 inst_cell_3_100 ( BL100, BLN100, WL3);
sram_cell_6t_3 inst_cell_2_100 ( BL100, BLN100, WL2);
sram_cell_6t_3 inst_cell_1_100 ( BL100, BLN100, WL1);
sram_cell_6t_3 inst_cell_0_100 ( BL100, BLN100, WL0);
sram_cell_6t_3 inst_cell_13_99 ( BL99, BLN99, WL13);
sram_cell_6t_3 inst_cell_12_99 ( BL99, BLN99, WL12);
sram_cell_6t_3 inst_cell_11_99 ( BL99, BLN99, WL11);
sram_cell_6t_3 inst_cell_10_99 ( BL99, BLN99, WL10);
sram_cell_6t_3 inst_cell_9_99 ( BL99, BLN99, WL9);
sram_cell_6t_3 inst_cell_8_99 ( BL99, BLN99, WL8);
sram_cell_6t_3 inst_cell_7_99 ( BL99, BLN99, WL7);
sram_cell_6t_3 inst_cell_6_99 ( BL99, BLN99, WL6);
sram_cell_6t_3 inst_cell_5_99 ( BL99, BLN99, WL5);
sram_cell_6t_3 inst_cell_4_99 ( BL99, BLN99, WL4);
sram_cell_6t_3 inst_cell_3_99 ( BL99, BLN99, WL3);
sram_cell_6t_3 inst_cell_2_99 ( BL99, BLN99, WL2);
sram_cell_6t_3 inst_cell_1_99 ( BL99, BLN99, WL1);
sram_cell_6t_3 inst_cell_0_99 ( BL99, BLN99, WL0);
sram_cell_6t_3 inst_cell_13_98 ( BL98, BLN98, WL13);
sram_cell_6t_3 inst_cell_12_98 ( BL98, BLN98, WL12);
sram_cell_6t_3 inst_cell_11_98 ( BL98, BLN98, WL11);
sram_cell_6t_3 inst_cell_10_98 ( BL98, BLN98, WL10);
sram_cell_6t_3 inst_cell_9_98 ( BL98, BLN98, WL9);
sram_cell_6t_3 inst_cell_8_98 ( BL98, BLN98, WL8);
sram_cell_6t_3 inst_cell_7_98 ( BL98, BLN98, WL7);
sram_cell_6t_3 inst_cell_6_98 ( BL98, BLN98, WL6);
sram_cell_6t_3 inst_cell_5_98 ( BL98, BLN98, WL5);
sram_cell_6t_3 inst_cell_4_98 ( BL98, BLN98, WL4);
sram_cell_6t_3 inst_cell_3_98 ( BL98, BLN98, WL3);
sram_cell_6t_3 inst_cell_2_98 ( BL98, BLN98, WL2);
sram_cell_6t_3 inst_cell_1_98 ( BL98, BLN98, WL1);
sram_cell_6t_3 inst_cell_0_98 ( BL98, BLN98, WL0);
sram_cell_6t_3 inst_cell_13_97 ( BL97, BLN97, WL13);
sram_cell_6t_3 inst_cell_12_97 ( BL97, BLN97, WL12);
sram_cell_6t_3 inst_cell_11_97 ( BL97, BLN97, WL11);
sram_cell_6t_3 inst_cell_10_97 ( BL97, BLN97, WL10);
sram_cell_6t_3 inst_cell_9_97 ( BL97, BLN97, WL9);
sram_cell_6t_3 inst_cell_8_97 ( BL97, BLN97, WL8);
sram_cell_6t_3 inst_cell_7_97 ( BL97, BLN97, WL7);
sram_cell_6t_3 inst_cell_6_97 ( BL97, BLN97, WL6);
sram_cell_6t_3 inst_cell_5_97 ( BL97, BLN97, WL5);
sram_cell_6t_3 inst_cell_4_97 ( BL97, BLN97, WL4);
sram_cell_6t_3 inst_cell_3_97 ( BL97, BLN97, WL3);
sram_cell_6t_3 inst_cell_2_97 ( BL97, BLN97, WL2);
sram_cell_6t_3 inst_cell_1_97 ( BL97, BLN97, WL1);
sram_cell_6t_3 inst_cell_0_97 ( BL97, BLN97, WL0);
sram_cell_6t_3 inst_cell_13_96 ( BL96, BLN96, WL13);
sram_cell_6t_3 inst_cell_12_96 ( BL96, BLN96, WL12);
sram_cell_6t_3 inst_cell_11_96 ( BL96, BLN96, WL11);
sram_cell_6t_3 inst_cell_10_96 ( BL96, BLN96, WL10);
sram_cell_6t_3 inst_cell_9_96 ( BL96, BLN96, WL9);
sram_cell_6t_3 inst_cell_8_96 ( BL96, BLN96, WL8);
sram_cell_6t_3 inst_cell_7_96 ( BL96, BLN96, WL7);
sram_cell_6t_3 inst_cell_6_96 ( BL96, BLN96, WL6);
sram_cell_6t_3 inst_cell_5_96 ( BL96, BLN96, WL5);
sram_cell_6t_3 inst_cell_4_96 ( BL96, BLN96, WL4);
sram_cell_6t_3 inst_cell_3_96 ( BL96, BLN96, WL3);
sram_cell_6t_3 inst_cell_2_96 ( BL96, BLN96, WL2);
sram_cell_6t_3 inst_cell_1_96 ( BL96, BLN96, WL1);
sram_cell_6t_3 inst_cell_0_96 ( BL96, BLN96, WL0);
sram_cell_6t_3 inst_cell_13_95 ( BL95, BLN95, WL13);
sram_cell_6t_3 inst_cell_12_95 ( BL95, BLN95, WL12);
sram_cell_6t_3 inst_cell_11_95 ( BL95, BLN95, WL11);
sram_cell_6t_3 inst_cell_10_95 ( BL95, BLN95, WL10);
sram_cell_6t_3 inst_cell_9_95 ( BL95, BLN95, WL9);
sram_cell_6t_3 inst_cell_8_95 ( BL95, BLN95, WL8);
sram_cell_6t_3 inst_cell_7_95 ( BL95, BLN95, WL7);
sram_cell_6t_3 inst_cell_6_95 ( BL95, BLN95, WL6);
sram_cell_6t_3 inst_cell_13_94 ( BL94, BLN94, WL13);
sram_cell_6t_3 inst_cell_12_94 ( BL94, BLN94, WL12);
sram_cell_6t_3 inst_cell_11_94 ( BL94, BLN94, WL11);
sram_cell_6t_3 inst_cell_10_94 ( BL94, BLN94, WL10);
sram_cell_6t_3 inst_cell_9_94 ( BL94, BLN94, WL9);
sram_cell_6t_3 inst_cell_8_94 ( BL94, BLN94, WL8);
sram_cell_6t_3 inst_cell_7_94 ( BL94, BLN94, WL7);
sram_cell_6t_3 inst_cell_6_94 ( BL94, BLN94, WL6);
sram_cell_6t_3 inst_cell_5_94 ( BL94, BLN94, WL5);
sram_cell_6t_3 inst_cell_4_94 ( BL94, BLN94, WL4);
sram_cell_6t_3 inst_cell_3_94 ( BL94, BLN94, WL3);
sram_cell_6t_3 inst_cell_2_94 ( BL94, BLN94, WL2);
sram_cell_6t_3 inst_cell_1_94 ( BL94, BLN94, WL1);
sram_cell_6t_3 inst_cell_0_94 ( BL94, BLN94, WL0);
sram_cell_6t_3 inst_cell_13_93 ( BL93, BLN93, WL13);
sram_cell_6t_3 inst_cell_12_93 ( BL93, BLN93, WL12);
sram_cell_6t_3 inst_cell_11_93 ( BL93, BLN93, WL11);
sram_cell_6t_3 inst_cell_10_93 ( BL93, BLN93, WL10);
sram_cell_6t_3 inst_cell_9_93 ( BL93, BLN93, WL9);
sram_cell_6t_3 inst_cell_8_93 ( BL93, BLN93, WL8);
sram_cell_6t_3 inst_cell_7_93 ( BL93, BLN93, WL7);
sram_cell_6t_3 inst_cell_6_93 ( BL93, BLN93, WL6);
sram_cell_6t_3 inst_cell_5_93 ( BL93, BLN93, WL5);
sram_cell_6t_3 inst_cell_4_93 ( BL93, BLN93, WL4);
sram_cell_6t_3 inst_cell_3_93 ( BL93, BLN93, WL3);
sram_cell_6t_3 inst_cell_2_93 ( BL93, BLN93, WL2);
sram_cell_6t_3 inst_cell_1_93 ( BL93, BLN93, WL1);
sram_cell_6t_3 inst_cell_0_93 ( BL93, BLN93, WL0);
sram_cell_6t_3 inst_cell_13_92 ( BL92, BLN92, WL13);
sram_cell_6t_3 inst_cell_12_92 ( BL92, BLN92, WL12);
sram_cell_6t_3 inst_cell_11_92 ( BL92, BLN92, WL11);
sram_cell_6t_3 inst_cell_10_92 ( BL92, BLN92, WL10);
sram_cell_6t_3 inst_cell_9_92 ( BL92, BLN92, WL9);
sram_cell_6t_3 inst_cell_8_92 ( BL92, BLN92, WL8);
sram_cell_6t_3 inst_cell_7_92 ( BL92, BLN92, WL7);
sram_cell_6t_3 inst_cell_6_92 ( BL92, BLN92, WL6);
sram_cell_6t_3 inst_cell_5_92 ( BL92, BLN92, WL5);
sram_cell_6t_3 inst_cell_4_92 ( BL92, BLN92, WL4);
sram_cell_6t_3 inst_cell_3_92 ( BL92, BLN92, WL3);
sram_cell_6t_3 inst_cell_2_92 ( BL92, BLN92, WL2);
sram_cell_6t_3 inst_cell_1_92 ( BL92, BLN92, WL1);
sram_cell_6t_3 inst_cell_0_92 ( BL92, BLN92, WL0);
sram_cell_6t_3 inst_cell_13_91 ( BL91, BLN91, WL13);
sram_cell_6t_3 inst_cell_12_91 ( BL91, BLN91, WL12);
sram_cell_6t_3 inst_cell_11_91 ( BL91, BLN91, WL11);
sram_cell_6t_3 inst_cell_10_91 ( BL91, BLN91, WL10);
sram_cell_6t_3 inst_cell_9_91 ( BL91, BLN91, WL9);
sram_cell_6t_3 inst_cell_8_91 ( BL91, BLN91, WL8);
sram_cell_6t_3 inst_cell_7_91 ( BL91, BLN91, WL7);
sram_cell_6t_3 inst_cell_6_91 ( BL91, BLN91, WL6);
sram_cell_6t_3 inst_cell_5_91 ( BL91, BLN91, WL5);
sram_cell_6t_3 inst_cell_4_91 ( BL91, BLN91, WL4);
sram_cell_6t_3 inst_cell_3_91 ( BL91, BLN91, WL3);
sram_cell_6t_3 inst_cell_2_91 ( BL91, BLN91, WL2);
sram_cell_6t_3 inst_cell_1_91 ( BL91, BLN91, WL1);
sram_cell_6t_3 inst_cell_0_91 ( BL91, BLN91, WL0);
sram_cell_6t_3 inst_cell_13_90 ( BL90, BLN90, WL13);
sram_cell_6t_3 inst_cell_12_90 ( BL90, BLN90, WL12);
sram_cell_6t_3 inst_cell_11_90 ( BL90, BLN90, WL11);
sram_cell_6t_3 inst_cell_10_90 ( BL90, BLN90, WL10);
sram_cell_6t_3 inst_cell_9_90 ( BL90, BLN90, WL9);
sram_cell_6t_3 inst_cell_8_90 ( BL90, BLN90, WL8);
sram_cell_6t_3 inst_cell_7_90 ( BL90, BLN90, WL7);
sram_cell_6t_3 inst_cell_6_90 ( BL90, BLN90, WL6);
sram_cell_6t_3 inst_cell_5_90 ( BL90, BLN90, WL5);
sram_cell_6t_3 inst_cell_4_90 ( BL90, BLN90, WL4);
sram_cell_6t_3 inst_cell_3_90 ( BL90, BLN90, WL3);
sram_cell_6t_3 inst_cell_2_90 ( BL90, BLN90, WL2);
sram_cell_6t_3 inst_cell_1_90 ( BL90, BLN90, WL1);
sram_cell_6t_3 inst_cell_0_90 ( BL90, BLN90, WL0);
sram_cell_6t_3 inst_cell_13_89 ( BL89, BLN89, WL13);
sram_cell_6t_3 inst_cell_12_89 ( BL89, BLN89, WL12);
sram_cell_6t_3 inst_cell_11_89 ( BL89, BLN89, WL11);
sram_cell_6t_3 inst_cell_10_89 ( BL89, BLN89, WL10);
sram_cell_6t_3 inst_cell_9_89 ( BL89, BLN89, WL9);
sram_cell_6t_3 inst_cell_8_89 ( BL89, BLN89, WL8);
sram_cell_6t_3 inst_cell_7_89 ( BL89, BLN89, WL7);
sram_cell_6t_3 inst_cell_6_89 ( BL89, BLN89, WL6);
sram_cell_6t_3 inst_cell_5_89 ( BL89, BLN89, WL5);
sram_cell_6t_3 inst_cell_4_89 ( BL89, BLN89, WL4);
sram_cell_6t_3 inst_cell_3_89 ( BL89, BLN89, WL3);
sram_cell_6t_3 inst_cell_2_89 ( BL89, BLN89, WL2);
sram_cell_6t_3 inst_cell_1_89 ( BL89, BLN89, WL1);
sram_cell_6t_3 inst_cell_0_89 ( BL89, BLN89, WL0);
sram_cell_6t_3 inst_cell_13_88 ( BL88, BLN88, WL13);
sram_cell_6t_3 inst_cell_12_88 ( BL88, BLN88, WL12);
sram_cell_6t_3 inst_cell_11_88 ( BL88, BLN88, WL11);
sram_cell_6t_3 inst_cell_10_88 ( BL88, BLN88, WL10);
sram_cell_6t_3 inst_cell_9_88 ( BL88, BLN88, WL9);
sram_cell_6t_3 inst_cell_8_88 ( BL88, BLN88, WL8);
sram_cell_6t_3 inst_cell_7_88 ( BL88, BLN88, WL7);
sram_cell_6t_3 inst_cell_6_88 ( BL88, BLN88, WL6);
sram_cell_6t_3 inst_cell_5_88 ( BL88, BLN88, WL5);
sram_cell_6t_3 inst_cell_4_88 ( BL88, BLN88, WL4);
sram_cell_6t_3 inst_cell_3_88 ( BL88, BLN88, WL3);
sram_cell_6t_3 inst_cell_2_88 ( BL88, BLN88, WL2);
sram_cell_6t_3 inst_cell_1_88 ( BL88, BLN88, WL1);
sram_cell_6t_3 inst_cell_0_88 ( BL88, BLN88, WL0);
sram_cell_6t_3 inst_cell_13_87 ( BL87, BLN87, WL13);
sram_cell_6t_3 inst_cell_12_87 ( BL87, BLN87, WL12);
sram_cell_6t_3 inst_cell_11_87 ( BL87, BLN87, WL11);
sram_cell_6t_3 inst_cell_10_87 ( BL87, BLN87, WL10);
sram_cell_6t_3 inst_cell_9_87 ( BL87, BLN87, WL9);
sram_cell_6t_3 inst_cell_8_87 ( BL87, BLN87, WL8);
sram_cell_6t_3 inst_cell_7_87 ( BL87, BLN87, WL7);
sram_cell_6t_3 inst_cell_6_87 ( BL87, BLN87, WL6);
sram_cell_6t_3 inst_cell_5_87 ( BL87, BLN87, WL5);
sram_cell_6t_3 inst_cell_4_87 ( BL87, BLN87, WL4);
sram_cell_6t_3 inst_cell_3_87 ( BL87, BLN87, WL3);
sram_cell_6t_3 inst_cell_2_87 ( BL87, BLN87, WL2);
sram_cell_6t_3 inst_cell_1_87 ( BL87, BLN87, WL1);
sram_cell_6t_3 inst_cell_0_87 ( BL87, BLN87, WL0);
sram_cell_6t_3 inst_cell_13_86 ( BL86, BLN86, WL13);
sram_cell_6t_3 inst_cell_12_86 ( BL86, BLN86, WL12);
sram_cell_6t_3 inst_cell_11_86 ( BL86, BLN86, WL11);
sram_cell_6t_3 inst_cell_10_86 ( BL86, BLN86, WL10);
sram_cell_6t_3 inst_cell_9_86 ( BL86, BLN86, WL9);
sram_cell_6t_3 inst_cell_8_86 ( BL86, BLN86, WL8);
sram_cell_6t_3 inst_cell_7_86 ( BL86, BLN86, WL7);
sram_cell_6t_3 inst_cell_6_86 ( BL86, BLN86, WL6);
sram_cell_6t_3 inst_cell_5_86 ( BL86, BLN86, WL5);
sram_cell_6t_3 inst_cell_4_86 ( BL86, BLN86, WL4);
sram_cell_6t_3 inst_cell_3_86 ( BL86, BLN86, WL3);
sram_cell_6t_3 inst_cell_2_86 ( BL86, BLN86, WL2);
sram_cell_6t_3 inst_cell_1_86 ( BL86, BLN86, WL1);
sram_cell_6t_3 inst_cell_0_86 ( BL86, BLN86, WL0);
sram_cell_6t_3 inst_cell_13_85 ( BL85, BLN85, WL13);
sram_cell_6t_3 inst_cell_12_85 ( BL85, BLN85, WL12);
sram_cell_6t_3 inst_cell_11_85 ( BL85, BLN85, WL11);
sram_cell_6t_3 inst_cell_10_85 ( BL85, BLN85, WL10);
sram_cell_6t_3 inst_cell_9_85 ( BL85, BLN85, WL9);
sram_cell_6t_3 inst_cell_8_85 ( BL85, BLN85, WL8);
sram_cell_6t_3 inst_cell_7_85 ( BL85, BLN85, WL7);
sram_cell_6t_3 inst_cell_6_85 ( BL85, BLN85, WL6);
sram_cell_6t_3 inst_cell_5_85 ( BL85, BLN85, WL5);
sram_cell_6t_3 inst_cell_4_85 ( BL85, BLN85, WL4);
sram_cell_6t_3 inst_cell_3_85 ( BL85, BLN85, WL3);
sram_cell_6t_3 inst_cell_2_85 ( BL85, BLN85, WL2);
sram_cell_6t_3 inst_cell_1_85 ( BL85, BLN85, WL1);
sram_cell_6t_3 inst_cell_0_85 ( BL85, BLN85, WL0);
sram_cell_6t_3 inst_cell_13_84 ( BL84, BLN84, WL13);
sram_cell_6t_3 inst_cell_12_84 ( BL84, BLN84, WL12);
sram_cell_6t_3 inst_cell_11_84 ( BL84, BLN84, WL11);
sram_cell_6t_3 inst_cell_10_84 ( BL84, BLN84, WL10);
sram_cell_6t_3 inst_cell_9_84 ( BL84, BLN84, WL9);
sram_cell_6t_3 inst_cell_8_84 ( BL84, BLN84, WL8);
sram_cell_6t_3 inst_cell_7_84 ( BL84, BLN84, WL7);
sram_cell_6t_3 inst_cell_6_84 ( BL84, BLN84, WL6);
sram_cell_6t_3 inst_cell_5_84 ( BL84, BLN84, WL5);
sram_cell_6t_3 inst_cell_4_84 ( BL84, BLN84, WL4);
sram_cell_6t_3 inst_cell_3_84 ( BL84, BLN84, WL3);
sram_cell_6t_3 inst_cell_2_84 ( BL84, BLN84, WL2);
sram_cell_6t_3 inst_cell_1_84 ( BL84, BLN84, WL1);
sram_cell_6t_3 inst_cell_0_84 ( BL84, BLN84, WL0);
sram_cell_6t_3 inst_cell_13_83 ( BL83, BLN83, WL13);
sram_cell_6t_3 inst_cell_12_83 ( BL83, BLN83, WL12);
sram_cell_6t_3 inst_cell_11_83 ( BL83, BLN83, WL11);
sram_cell_6t_3 inst_cell_10_83 ( BL83, BLN83, WL10);
sram_cell_6t_3 inst_cell_9_83 ( BL83, BLN83, WL9);
sram_cell_6t_3 inst_cell_8_83 ( BL83, BLN83, WL8);
sram_cell_6t_3 inst_cell_7_83 ( BL83, BLN83, WL7);
sram_cell_6t_3 inst_cell_6_83 ( BL83, BLN83, WL6);
sram_cell_6t_3 inst_cell_5_83 ( BL83, BLN83, WL5);
sram_cell_6t_3 inst_cell_4_83 ( BL83, BLN83, WL4);
sram_cell_6t_3 inst_cell_3_83 ( BL83, BLN83, WL3);
sram_cell_6t_3 inst_cell_2_83 ( BL83, BLN83, WL2);
sram_cell_6t_3 inst_cell_1_83 ( BL83, BLN83, WL1);
sram_cell_6t_3 inst_cell_0_83 ( BL83, BLN83, WL0);
sram_cell_6t_3 inst_cell_13_82 ( BL82, BLN82, WL13);
sram_cell_6t_3 inst_cell_12_82 ( BL82, BLN82, WL12);
sram_cell_6t_3 inst_cell_11_82 ( BL82, BLN82, WL11);
sram_cell_6t_3 inst_cell_10_82 ( BL82, BLN82, WL10);
sram_cell_6t_3 inst_cell_9_82 ( BL82, BLN82, WL9);
sram_cell_6t_3 inst_cell_8_82 ( BL82, BLN82, WL8);
sram_cell_6t_3 inst_cell_7_82 ( BL82, BLN82, WL7);
sram_cell_6t_3 inst_cell_6_82 ( BL82, BLN82, WL6);
sram_cell_6t_3 inst_cell_5_82 ( BL82, BLN82, WL5);
sram_cell_6t_3 inst_cell_4_82 ( BL82, BLN82, WL4);
sram_cell_6t_3 inst_cell_3_82 ( BL82, BLN82, WL3);
sram_cell_6t_3 inst_cell_2_82 ( BL82, BLN82, WL2);
sram_cell_6t_3 inst_cell_1_82 ( BL82, BLN82, WL1);
sram_cell_6t_3 inst_cell_0_82 ( BL82, BLN82, WL0);
sram_cell_6t_3 inst_cell_13_81 ( BL81, BLN81, WL13);
sram_cell_6t_3 inst_cell_12_81 ( BL81, BLN81, WL12);
sram_cell_6t_3 inst_cell_11_81 ( BL81, BLN81, WL11);
sram_cell_6t_3 inst_cell_10_81 ( BL81, BLN81, WL10);
sram_cell_6t_3 inst_cell_9_81 ( BL81, BLN81, WL9);
sram_cell_6t_3 inst_cell_8_81 ( BL81, BLN81, WL8);
sram_cell_6t_3 inst_cell_7_81 ( BL81, BLN81, WL7);
sram_cell_6t_3 inst_cell_6_81 ( BL81, BLN81, WL6);
sram_cell_6t_3 inst_cell_5_81 ( BL81, BLN81, WL5);
sram_cell_6t_3 inst_cell_4_81 ( BL81, BLN81, WL4);
sram_cell_6t_3 inst_cell_3_81 ( BL81, BLN81, WL3);
sram_cell_6t_3 inst_cell_2_81 ( BL81, BLN81, WL2);
sram_cell_6t_3 inst_cell_1_81 ( BL81, BLN81, WL1);
sram_cell_6t_3 inst_cell_0_81 ( BL81, BLN81, WL0);
sram_cell_6t_3 inst_cell_13_80 ( BL80, BLN80, WL13);
sram_cell_6t_3 inst_cell_12_80 ( BL80, BLN80, WL12);
sram_cell_6t_3 inst_cell_11_80 ( BL80, BLN80, WL11);
sram_cell_6t_3 inst_cell_10_80 ( BL80, BLN80, WL10);
sram_cell_6t_3 inst_cell_9_80 ( BL80, BLN80, WL9);
sram_cell_6t_3 inst_cell_8_80 ( BL80, BLN80, WL8);
sram_cell_6t_3 inst_cell_7_80 ( BL80, BLN80, WL7);
sram_cell_6t_3 inst_cell_6_80 ( BL80, BLN80, WL6);
sram_cell_6t_3 inst_cell_5_80 ( BL80, BLN80, WL5);
sram_cell_6t_3 inst_cell_4_80 ( BL80, BLN80, WL4);
sram_cell_6t_3 inst_cell_3_80 ( BL80, BLN80, WL3);
sram_cell_6t_3 inst_cell_2_80 ( BL80, BLN80, WL2);
sram_cell_6t_3 inst_cell_1_80 ( BL80, BLN80, WL1);
sram_cell_6t_3 inst_cell_0_80 ( BL80, BLN80, WL0);
sram_cell_6t_3 inst_cell_13_79 ( BL79, BLN79, WL13);
sram_cell_6t_3 inst_cell_12_79 ( BL79, BLN79, WL12);
sram_cell_6t_3 inst_cell_11_79 ( BL79, BLN79, WL11);
sram_cell_6t_3 inst_cell_10_79 ( BL79, BLN79, WL10);
sram_cell_6t_3 inst_cell_9_79 ( BL79, BLN79, WL9);
sram_cell_6t_3 inst_cell_8_79 ( BL79, BLN79, WL8);
sram_cell_6t_3 inst_cell_7_79 ( BL79, BLN79, WL7);
sram_cell_6t_3 inst_cell_6_79 ( BL79, BLN79, WL6);
sram_cell_6t_3 inst_cell_5_79 ( BL79, BLN79, WL5);
sram_cell_6t_3 inst_cell_4_79 ( BL79, BLN79, WL4);
sram_cell_6t_3 inst_cell_3_79 ( BL79, BLN79, WL3);
sram_cell_6t_3 inst_cell_2_79 ( BL79, BLN79, WL2);
sram_cell_6t_3 inst_cell_1_79 ( BL79, BLN79, WL1);
sram_cell_6t_3 inst_cell_0_79 ( BL79, BLN79, WL0);
sram_cell_6t_3 inst_cell_13_78 ( BL78, BLN78, WL13);
sram_cell_6t_3 inst_cell_12_78 ( BL78, BLN78, WL12);
sram_cell_6t_3 inst_cell_11_78 ( BL78, BLN78, WL11);
sram_cell_6t_3 inst_cell_10_78 ( BL78, BLN78, WL10);
sram_cell_6t_3 inst_cell_9_78 ( BL78, BLN78, WL9);
sram_cell_6t_3 inst_cell_8_78 ( BL78, BLN78, WL8);
sram_cell_6t_3 inst_cell_7_78 ( BL78, BLN78, WL7);
sram_cell_6t_3 inst_cell_6_78 ( BL78, BLN78, WL6);
sram_cell_6t_3 inst_cell_5_78 ( BL78, BLN78, WL5);
sram_cell_6t_3 inst_cell_4_78 ( BL78, BLN78, WL4);
sram_cell_6t_3 inst_cell_3_78 ( BL78, BLN78, WL3);
sram_cell_6t_3 inst_cell_2_78 ( BL78, BLN78, WL2);
sram_cell_6t_3 inst_cell_1_78 ( BL78, BLN78, WL1);
sram_cell_6t_3 inst_cell_0_78 ( BL78, BLN78, WL0);
sram_cell_6t_3 inst_cell_13_77 ( BL77, BLN77, WL13);
sram_cell_6t_3 inst_cell_12_77 ( BL77, BLN77, WL12);
sram_cell_6t_3 inst_cell_11_77 ( BL77, BLN77, WL11);
sram_cell_6t_3 inst_cell_10_77 ( BL77, BLN77, WL10);
sram_cell_6t_3 inst_cell_9_77 ( BL77, BLN77, WL9);
sram_cell_6t_3 inst_cell_8_77 ( BL77, BLN77, WL8);
sram_cell_6t_3 inst_cell_7_77 ( BL77, BLN77, WL7);
sram_cell_6t_3 inst_cell_6_77 ( BL77, BLN77, WL6);
sram_cell_6t_3 inst_cell_5_77 ( BL77, BLN77, WL5);
sram_cell_6t_3 inst_cell_4_77 ( BL77, BLN77, WL4);
sram_cell_6t_3 inst_cell_3_77 ( BL77, BLN77, WL3);
sram_cell_6t_3 inst_cell_2_77 ( BL77, BLN77, WL2);
sram_cell_6t_3 inst_cell_1_77 ( BL77, BLN77, WL1);
sram_cell_6t_3 inst_cell_0_77 ( BL77, BLN77, WL0);
sram_cell_6t_3 inst_cell_13_76 ( BL76, BLN76, WL13);
sram_cell_6t_3 inst_cell_12_76 ( BL76, BLN76, WL12);
sram_cell_6t_3 inst_cell_11_76 ( BL76, BLN76, WL11);
sram_cell_6t_3 inst_cell_10_76 ( BL76, BLN76, WL10);
sram_cell_6t_3 inst_cell_9_76 ( BL76, BLN76, WL9);
sram_cell_6t_3 inst_cell_8_76 ( BL76, BLN76, WL8);
sram_cell_6t_3 inst_cell_7_76 ( BL76, BLN76, WL7);
sram_cell_6t_3 inst_cell_6_76 ( BL76, BLN76, WL6);
sram_cell_6t_3 inst_cell_5_76 ( BL76, BLN76, WL5);
sram_cell_6t_3 inst_cell_4_76 ( BL76, BLN76, WL4);
sram_cell_6t_3 inst_cell_3_76 ( BL76, BLN76, WL3);
sram_cell_6t_3 inst_cell_2_76 ( BL76, BLN76, WL2);
sram_cell_6t_3 inst_cell_1_76 ( BL76, BLN76, WL1);
sram_cell_6t_3 inst_cell_0_76 ( BL76, BLN76, WL0);
sram_cell_6t_3 inst_cell_13_75 ( BL75, BLN75, WL13);
sram_cell_6t_3 inst_cell_12_75 ( BL75, BLN75, WL12);
sram_cell_6t_3 inst_cell_11_75 ( BL75, BLN75, WL11);
sram_cell_6t_3 inst_cell_10_75 ( BL75, BLN75, WL10);
sram_cell_6t_3 inst_cell_9_75 ( BL75, BLN75, WL9);
sram_cell_6t_3 inst_cell_8_75 ( BL75, BLN75, WL8);
sram_cell_6t_3 inst_cell_7_75 ( BL75, BLN75, WL7);
sram_cell_6t_3 inst_cell_6_75 ( BL75, BLN75, WL6);
sram_cell_6t_3 inst_cell_5_75 ( BL75, BLN75, WL5);
sram_cell_6t_3 inst_cell_4_75 ( BL75, BLN75, WL4);
sram_cell_6t_3 inst_cell_3_75 ( BL75, BLN75, WL3);
sram_cell_6t_3 inst_cell_2_75 ( BL75, BLN75, WL2);
sram_cell_6t_3 inst_cell_1_75 ( BL75, BLN75, WL1);
sram_cell_6t_3 inst_cell_0_75 ( BL75, BLN75, WL0);
sram_cell_6t_3 inst_cell_13_74 ( BL74, BLN74, WL13);
sram_cell_6t_3 inst_cell_12_74 ( BL74, BLN74, WL12);
sram_cell_6t_3 inst_cell_11_74 ( BL74, BLN74, WL11);
sram_cell_6t_3 inst_cell_10_74 ( BL74, BLN74, WL10);
sram_cell_6t_3 inst_cell_9_74 ( BL74, BLN74, WL9);
sram_cell_6t_3 inst_cell_8_74 ( BL74, BLN74, WL8);
sram_cell_6t_3 inst_cell_7_74 ( BL74, BLN74, WL7);
sram_cell_6t_3 inst_cell_6_74 ( BL74, BLN74, WL6);
sram_cell_6t_3 inst_cell_5_74 ( BL74, BLN74, WL5);
sram_cell_6t_3 inst_cell_4_74 ( BL74, BLN74, WL4);
sram_cell_6t_3 inst_cell_3_74 ( BL74, BLN74, WL3);
sram_cell_6t_3 inst_cell_2_74 ( BL74, BLN74, WL2);
sram_cell_6t_3 inst_cell_1_74 ( BL74, BLN74, WL1);
sram_cell_6t_3 inst_cell_0_74 ( BL74, BLN74, WL0);
sram_cell_6t_3 inst_cell_13_73 ( BL73, BLN73, WL13);
sram_cell_6t_3 inst_cell_12_73 ( BL73, BLN73, WL12);
sram_cell_6t_3 inst_cell_11_73 ( BL73, BLN73, WL11);
sram_cell_6t_3 inst_cell_10_73 ( BL73, BLN73, WL10);
sram_cell_6t_3 inst_cell_9_73 ( BL73, BLN73, WL9);
sram_cell_6t_3 inst_cell_8_73 ( BL73, BLN73, WL8);
sram_cell_6t_3 inst_cell_7_73 ( BL73, BLN73, WL7);
sram_cell_6t_3 inst_cell_6_73 ( BL73, BLN73, WL6);
sram_cell_6t_3 inst_cell_5_73 ( BL73, BLN73, WL5);
sram_cell_6t_3 inst_cell_4_73 ( BL73, BLN73, WL4);
sram_cell_6t_3 inst_cell_3_73 ( BL73, BLN73, WL3);
sram_cell_6t_3 inst_cell_2_73 ( BL73, BLN73, WL2);
sram_cell_6t_3 inst_cell_1_73 ( BL73, BLN73, WL1);
sram_cell_6t_3 inst_cell_0_73 ( BL73, BLN73, WL0);
sram_cell_6t_3 inst_cell_13_72 ( BL72, BLN72, WL13);
sram_cell_6t_3 inst_cell_12_72 ( BL72, BLN72, WL12);
sram_cell_6t_3 inst_cell_11_72 ( BL72, BLN72, WL11);
sram_cell_6t_3 inst_cell_10_72 ( BL72, BLN72, WL10);
sram_cell_6t_3 inst_cell_9_72 ( BL72, BLN72, WL9);
sram_cell_6t_3 inst_cell_8_72 ( BL72, BLN72, WL8);
sram_cell_6t_3 inst_cell_7_72 ( BL72, BLN72, WL7);
sram_cell_6t_3 inst_cell_6_72 ( BL72, BLN72, WL6);
sram_cell_6t_3 inst_cell_5_72 ( BL72, BLN72, WL5);
sram_cell_6t_3 inst_cell_4_72 ( BL72, BLN72, WL4);
sram_cell_6t_3 inst_cell_3_72 ( BL72, BLN72, WL3);
sram_cell_6t_3 inst_cell_2_72 ( BL72, BLN72, WL2);
sram_cell_6t_3 inst_cell_1_72 ( BL72, BLN72, WL1);
sram_cell_6t_3 inst_cell_0_72 ( BL72, BLN72, WL0);
sram_cell_6t_3 inst_cell_13_71 ( BL71, BLN71, WL13);
sram_cell_6t_3 inst_cell_12_71 ( BL71, BLN71, WL12);
sram_cell_6t_3 inst_cell_11_71 ( BL71, BLN71, WL11);
sram_cell_6t_3 inst_cell_10_71 ( BL71, BLN71, WL10);
sram_cell_6t_3 inst_cell_9_71 ( BL71, BLN71, WL9);
sram_cell_6t_3 inst_cell_8_71 ( BL71, BLN71, WL8);
sram_cell_6t_3 inst_cell_7_71 ( BL71, BLN71, WL7);
sram_cell_6t_3 inst_cell_6_71 ( BL71, BLN71, WL6);
sram_cell_6t_3 inst_cell_5_71 ( BL71, BLN71, WL5);
sram_cell_6t_3 inst_cell_4_71 ( BL71, BLN71, WL4);
sram_cell_6t_3 inst_cell_3_71 ( BL71, BLN71, WL3);
sram_cell_6t_3 inst_cell_2_71 ( BL71, BLN71, WL2);
sram_cell_6t_3 inst_cell_1_71 ( BL71, BLN71, WL1);
sram_cell_6t_3 inst_cell_0_71 ( BL71, BLN71, WL0);
sram_cell_6t_3 inst_cell_13_70 ( BL70, BLN70, WL13);
sram_cell_6t_3 inst_cell_12_70 ( BL70, BLN70, WL12);
sram_cell_6t_3 inst_cell_11_70 ( BL70, BLN70, WL11);
sram_cell_6t_3 inst_cell_10_70 ( BL70, BLN70, WL10);
sram_cell_6t_3 inst_cell_9_70 ( BL70, BLN70, WL9);
sram_cell_6t_3 inst_cell_8_70 ( BL70, BLN70, WL8);
sram_cell_6t_3 inst_cell_7_70 ( BL70, BLN70, WL7);
sram_cell_6t_3 inst_cell_6_70 ( BL70, BLN70, WL6);
sram_cell_6t_3 inst_cell_5_70 ( BL70, BLN70, WL5);
sram_cell_6t_3 inst_cell_4_70 ( BL70, BLN70, WL4);
sram_cell_6t_3 inst_cell_3_70 ( BL70, BLN70, WL3);
sram_cell_6t_3 inst_cell_2_70 ( BL70, BLN70, WL2);
sram_cell_6t_3 inst_cell_1_70 ( BL70, BLN70, WL1);
sram_cell_6t_3 inst_cell_0_70 ( BL70, BLN70, WL0);
sram_cell_6t_3 inst_cell_13_69 ( BL69, BLN69, WL13);
sram_cell_6t_3 inst_cell_12_69 ( BL69, BLN69, WL12);
sram_cell_6t_3 inst_cell_11_69 ( BL69, BLN69, WL11);
sram_cell_6t_3 inst_cell_10_69 ( BL69, BLN69, WL10);
sram_cell_6t_3 inst_cell_9_69 ( BL69, BLN69, WL9);
sram_cell_6t_3 inst_cell_8_69 ( BL69, BLN69, WL8);
sram_cell_6t_3 inst_cell_7_69 ( BL69, BLN69, WL7);
sram_cell_6t_3 inst_cell_6_69 ( BL69, BLN69, WL6);
sram_cell_6t_3 inst_cell_5_69 ( BL69, BLN69, WL5);
sram_cell_6t_3 inst_cell_4_69 ( BL69, BLN69, WL4);
sram_cell_6t_3 inst_cell_3_69 ( BL69, BLN69, WL3);
sram_cell_6t_3 inst_cell_2_69 ( BL69, BLN69, WL2);
sram_cell_6t_3 inst_cell_1_69 ( BL69, BLN69, WL1);
sram_cell_6t_3 inst_cell_0_69 ( BL69, BLN69, WL0);
sram_cell_6t_3 inst_cell_13_68 ( BL68, BLN68, WL13);
sram_cell_6t_3 inst_cell_12_68 ( BL68, BLN68, WL12);
sram_cell_6t_3 inst_cell_11_68 ( BL68, BLN68, WL11);
sram_cell_6t_3 inst_cell_10_68 ( BL68, BLN68, WL10);
sram_cell_6t_3 inst_cell_9_68 ( BL68, BLN68, WL9);
sram_cell_6t_3 inst_cell_8_68 ( BL68, BLN68, WL8);
sram_cell_6t_3 inst_cell_7_68 ( BL68, BLN68, WL7);
sram_cell_6t_3 inst_cell_6_68 ( BL68, BLN68, WL6);
sram_cell_6t_3 inst_cell_5_68 ( BL68, BLN68, WL5);
sram_cell_6t_3 inst_cell_4_68 ( BL68, BLN68, WL4);
sram_cell_6t_3 inst_cell_3_68 ( BL68, BLN68, WL3);
sram_cell_6t_3 inst_cell_2_68 ( BL68, BLN68, WL2);
sram_cell_6t_3 inst_cell_1_68 ( BL68, BLN68, WL1);
sram_cell_6t_3 inst_cell_0_68 ( BL68, BLN68, WL0);
sram_cell_6t_3 inst_cell_13_67 ( BL67, BLN67, WL13);
sram_cell_6t_3 inst_cell_12_67 ( BL67, BLN67, WL12);
sram_cell_6t_3 inst_cell_11_67 ( BL67, BLN67, WL11);
sram_cell_6t_3 inst_cell_10_67 ( BL67, BLN67, WL10);
sram_cell_6t_3 inst_cell_9_67 ( BL67, BLN67, WL9);
sram_cell_6t_3 inst_cell_8_67 ( BL67, BLN67, WL8);
sram_cell_6t_3 inst_cell_7_67 ( BL67, BLN67, WL7);
sram_cell_6t_3 inst_cell_6_67 ( BL67, BLN67, WL6);
sram_cell_6t_3 inst_cell_5_67 ( BL67, BLN67, WL5);
sram_cell_6t_3 inst_cell_4_67 ( BL67, BLN67, WL4);
sram_cell_6t_3 inst_cell_3_67 ( BL67, BLN67, WL3);
sram_cell_6t_3 inst_cell_2_67 ( BL67, BLN67, WL2);
sram_cell_6t_3 inst_cell_1_67 ( BL67, BLN67, WL1);
sram_cell_6t_3 inst_cell_0_67 ( BL67, BLN67, WL0);
sram_cell_6t_3 inst_cell_13_66 ( BL66, BLN66, WL13);
sram_cell_6t_3 inst_cell_12_66 ( BL66, BLN66, WL12);
sram_cell_6t_3 inst_cell_11_66 ( BL66, BLN66, WL11);
sram_cell_6t_3 inst_cell_10_66 ( BL66, BLN66, WL10);
sram_cell_6t_3 inst_cell_9_66 ( BL66, BLN66, WL9);
sram_cell_6t_3 inst_cell_8_66 ( BL66, BLN66, WL8);
sram_cell_6t_3 inst_cell_7_66 ( BL66, BLN66, WL7);
sram_cell_6t_3 inst_cell_6_66 ( BL66, BLN66, WL6);
sram_cell_6t_3 inst_cell_5_66 ( BL66, BLN66, WL5);
sram_cell_6t_3 inst_cell_4_66 ( BL66, BLN66, WL4);
sram_cell_6t_3 inst_cell_3_66 ( BL66, BLN66, WL3);
sram_cell_6t_3 inst_cell_2_66 ( BL66, BLN66, WL2);
sram_cell_6t_3 inst_cell_1_66 ( BL66, BLN66, WL1);
sram_cell_6t_3 inst_cell_0_66 ( BL66, BLN66, WL0);
sram_cell_6t_3 inst_cell_13_65 ( BL65, BLN65, WL13);
sram_cell_6t_3 inst_cell_12_65 ( BL65, BLN65, WL12);
sram_cell_6t_3 inst_cell_11_65 ( BL65, BLN65, WL11);
sram_cell_6t_3 inst_cell_10_65 ( BL65, BLN65, WL10);
sram_cell_6t_3 inst_cell_9_65 ( BL65, BLN65, WL9);
sram_cell_6t_3 inst_cell_8_65 ( BL65, BLN65, WL8);
sram_cell_6t_3 inst_cell_7_65 ( BL65, BLN65, WL7);
sram_cell_6t_3 inst_cell_6_65 ( BL65, BLN65, WL6);
sram_cell_6t_3 inst_cell_5_65 ( BL65, BLN65, WL5);
sram_cell_6t_3 inst_cell_4_65 ( BL65, BLN65, WL4);
sram_cell_6t_3 inst_cell_3_65 ( BL65, BLN65, WL3);
sram_cell_6t_3 inst_cell_2_65 ( BL65, BLN65, WL2);
sram_cell_6t_3 inst_cell_1_65 ( BL65, BLN65, WL1);
sram_cell_6t_3 inst_cell_0_65 ( BL65, BLN65, WL0);
sram_cell_6t_3 inst_cell_13_64 ( BL64, BLN64, WL13);
sram_cell_6t_3 inst_cell_12_64 ( BL64, BLN64, WL12);
sram_cell_6t_3 inst_cell_11_64 ( BL64, BLN64, WL11);
sram_cell_6t_3 inst_cell_10_64 ( BL64, BLN64, WL10);
sram_cell_6t_3 inst_cell_9_64 ( BL64, BLN64, WL9);
sram_cell_6t_3 inst_cell_8_64 ( BL64, BLN64, WL8);
sram_cell_6t_3 inst_cell_7_64 ( BL64, BLN64, WL7);
sram_cell_6t_3 inst_cell_6_64 ( BL64, BLN64, WL6);
sram_cell_6t_3 inst_cell_5_64 ( BL64, BLN64, WL5);
sram_cell_6t_3 inst_cell_4_64 ( BL64, BLN64, WL4);
sram_cell_6t_3 inst_cell_3_64 ( BL64, BLN64, WL3);
sram_cell_6t_3 inst_cell_2_64 ( BL64, BLN64, WL2);
sram_cell_6t_3 inst_cell_1_64 ( BL64, BLN64, WL1);
sram_cell_6t_3 inst_cell_0_64 ( BL64, BLN64, WL0);
sram_cell_6t_3 inst_cell_13_63 ( BL63, BLN63, WL13);
sram_cell_6t_3 inst_cell_12_63 ( BL63, BLN63, WL12);
sram_cell_6t_3 inst_cell_11_63 ( BL63, BLN63, WL11);
sram_cell_6t_3 inst_cell_10_63 ( BL63, BLN63, WL10);
sram_cell_6t_3 inst_cell_9_63 ( BL63, BLN63, WL9);
sram_cell_6t_3 inst_cell_8_63 ( BL63, BLN63, WL8);
sram_cell_6t_3 inst_cell_7_63 ( BL63, BLN63, WL7);
sram_cell_6t_3 inst_cell_6_63 ( BL63, BLN63, WL6);
sram_cell_6t_3 inst_cell_5_63 ( BL63, BLN63, WL5);
sram_cell_6t_3 inst_cell_4_63 ( BL63, BLN63, WL4);
sram_cell_6t_3 inst_cell_3_63 ( BL63, BLN63, WL3);
sram_cell_6t_3 inst_cell_2_63 ( BL63, BLN63, WL2);
sram_cell_6t_3 inst_cell_1_63 ( BL63, BLN63, WL1);
sram_cell_6t_3 inst_cell_0_63 ( BL63, BLN63, WL0);
sram_cell_6t_3 inst_cell_13_62 ( BL62, BLN62, WL13);
sram_cell_6t_3 inst_cell_12_62 ( BL62, BLN62, WL12);
sram_cell_6t_3 inst_cell_11_62 ( BL62, BLN62, WL11);
sram_cell_6t_3 inst_cell_10_62 ( BL62, BLN62, WL10);
sram_cell_6t_3 inst_cell_9_62 ( BL62, BLN62, WL9);
sram_cell_6t_3 inst_cell_8_62 ( BL62, BLN62, WL8);
sram_cell_6t_3 inst_cell_7_62 ( BL62, BLN62, WL7);
sram_cell_6t_3 inst_cell_6_62 ( BL62, BLN62, WL6);
sram_cell_6t_3 inst_cell_13_61 ( BL61, BLN61, WL13);
sram_cell_6t_3 inst_cell_12_61 ( BL61, BLN61, WL12);
sram_cell_6t_3 inst_cell_11_61 ( BL61, BLN61, WL11);
sram_cell_6t_3 inst_cell_10_61 ( BL61, BLN61, WL10);
sram_cell_6t_3 inst_cell_9_61 ( BL61, BLN61, WL9);
sram_cell_6t_3 inst_cell_8_61 ( BL61, BLN61, WL8);
sram_cell_6t_3 inst_cell_7_61 ( BL61, BLN61, WL7);
sram_cell_6t_3 inst_cell_6_61 ( BL61, BLN61, WL6);
sram_cell_6t_3 inst_cell_5_61 ( BL61, BLN61, WL5);
sram_cell_6t_3 inst_cell_4_61 ( BL61, BLN61, WL4);
sram_cell_6t_3 inst_cell_3_61 ( BL61, BLN61, WL3);
sram_cell_6t_3 inst_cell_2_61 ( BL61, BLN61, WL2);
sram_cell_6t_3 inst_cell_1_61 ( BL61, BLN61, WL1);
sram_cell_6t_3 inst_cell_0_61 ( BL61, BLN61, WL0);
sram_cell_6t_3 inst_cell_13_60 ( BL60, BLN60, WL13);
sram_cell_6t_3 inst_cell_12_60 ( BL60, BLN60, WL12);
sram_cell_6t_3 inst_cell_11_60 ( BL60, BLN60, WL11);
sram_cell_6t_3 inst_cell_10_60 ( BL60, BLN60, WL10);
sram_cell_6t_3 inst_cell_9_60 ( BL60, BLN60, WL9);
sram_cell_6t_3 inst_cell_8_60 ( BL60, BLN60, WL8);
sram_cell_6t_3 inst_cell_7_60 ( BL60, BLN60, WL7);
sram_cell_6t_3 inst_cell_6_60 ( BL60, BLN60, WL6);
sram_cell_6t_3 inst_cell_5_60 ( BL60, BLN60, WL5);
sram_cell_6t_3 inst_cell_4_60 ( BL60, BLN60, WL4);
sram_cell_6t_3 inst_cell_3_60 ( BL60, BLN60, WL3);
sram_cell_6t_3 inst_cell_2_60 ( BL60, BLN60, WL2);
sram_cell_6t_3 inst_cell_1_60 ( BL60, BLN60, WL1);
sram_cell_6t_3 inst_cell_0_60 ( BL60, BLN60, WL0);
sram_cell_6t_3 inst_cell_13_59 ( BL59, BLN59, WL13);
sram_cell_6t_3 inst_cell_12_59 ( BL59, BLN59, WL12);
sram_cell_6t_3 inst_cell_11_59 ( BL59, BLN59, WL11);
sram_cell_6t_3 inst_cell_10_59 ( BL59, BLN59, WL10);
sram_cell_6t_3 inst_cell_9_59 ( BL59, BLN59, WL9);
sram_cell_6t_3 inst_cell_8_59 ( BL59, BLN59, WL8);
sram_cell_6t_3 inst_cell_7_59 ( BL59, BLN59, WL7);
sram_cell_6t_3 inst_cell_6_59 ( BL59, BLN59, WL6);
sram_cell_6t_3 inst_cell_5_59 ( BL59, BLN59, WL5);
sram_cell_6t_3 inst_cell_4_59 ( BL59, BLN59, WL4);
sram_cell_6t_3 inst_cell_3_59 ( BL59, BLN59, WL3);
sram_cell_6t_3 inst_cell_2_59 ( BL59, BLN59, WL2);
sram_cell_6t_3 inst_cell_1_59 ( BL59, BLN59, WL1);
sram_cell_6t_3 inst_cell_0_59 ( BL59, BLN59, WL0);
sram_cell_6t_3 inst_cell_13_58 ( BL58, BLN58, WL13);
sram_cell_6t_3 inst_cell_12_58 ( BL58, BLN58, WL12);
sram_cell_6t_3 inst_cell_11_58 ( BL58, BLN58, WL11);
sram_cell_6t_3 inst_cell_10_58 ( BL58, BLN58, WL10);
sram_cell_6t_3 inst_cell_9_58 ( BL58, BLN58, WL9);
sram_cell_6t_3 inst_cell_8_58 ( BL58, BLN58, WL8);
sram_cell_6t_3 inst_cell_7_58 ( BL58, BLN58, WL7);
sram_cell_6t_3 inst_cell_6_58 ( BL58, BLN58, WL6);
sram_cell_6t_3 inst_cell_5_58 ( BL58, BLN58, WL5);
sram_cell_6t_3 inst_cell_4_58 ( BL58, BLN58, WL4);
sram_cell_6t_3 inst_cell_3_58 ( BL58, BLN58, WL3);
sram_cell_6t_3 inst_cell_2_58 ( BL58, BLN58, WL2);
sram_cell_6t_3 inst_cell_1_58 ( BL58, BLN58, WL1);
sram_cell_6t_3 inst_cell_0_58 ( BL58, BLN58, WL0);
sram_cell_6t_3 inst_cell_13_57 ( BL57, BLN57, WL13);
sram_cell_6t_3 inst_cell_12_57 ( BL57, BLN57, WL12);
sram_cell_6t_3 inst_cell_11_57 ( BL57, BLN57, WL11);
sram_cell_6t_3 inst_cell_10_57 ( BL57, BLN57, WL10);
sram_cell_6t_3 inst_cell_9_57 ( BL57, BLN57, WL9);
sram_cell_6t_3 inst_cell_8_57 ( BL57, BLN57, WL8);
sram_cell_6t_3 inst_cell_7_57 ( BL57, BLN57, WL7);
sram_cell_6t_3 inst_cell_6_57 ( BL57, BLN57, WL6);
sram_cell_6t_3 inst_cell_5_57 ( BL57, BLN57, WL5);
sram_cell_6t_3 inst_cell_4_57 ( BL57, BLN57, WL4);
sram_cell_6t_3 inst_cell_3_57 ( BL57, BLN57, WL3);
sram_cell_6t_3 inst_cell_2_57 ( BL57, BLN57, WL2);
sram_cell_6t_3 inst_cell_1_57 ( BL57, BLN57, WL1);
sram_cell_6t_3 inst_cell_0_57 ( BL57, BLN57, WL0);
sram_cell_6t_3 inst_cell_13_56 ( BL56, BLN56, WL13);
sram_cell_6t_3 inst_cell_12_56 ( BL56, BLN56, WL12);
sram_cell_6t_3 inst_cell_11_56 ( BL56, BLN56, WL11);
sram_cell_6t_3 inst_cell_10_56 ( BL56, BLN56, WL10);
sram_cell_6t_3 inst_cell_9_56 ( BL56, BLN56, WL9);
sram_cell_6t_3 inst_cell_8_56 ( BL56, BLN56, WL8);
sram_cell_6t_3 inst_cell_7_56 ( BL56, BLN56, WL7);
sram_cell_6t_3 inst_cell_6_56 ( BL56, BLN56, WL6);
sram_cell_6t_3 inst_cell_5_56 ( BL56, BLN56, WL5);
sram_cell_6t_3 inst_cell_4_56 ( BL56, BLN56, WL4);
sram_cell_6t_3 inst_cell_3_56 ( BL56, BLN56, WL3);
sram_cell_6t_3 inst_cell_2_56 ( BL56, BLN56, WL2);
sram_cell_6t_3 inst_cell_1_56 ( BL56, BLN56, WL1);
sram_cell_6t_3 inst_cell_0_56 ( BL56, BLN56, WL0);
sram_cell_6t_3 inst_cell_13_55 ( BL55, BLN55, WL13);
sram_cell_6t_3 inst_cell_12_55 ( BL55, BLN55, WL12);
sram_cell_6t_3 inst_cell_11_55 ( BL55, BLN55, WL11);
sram_cell_6t_3 inst_cell_10_55 ( BL55, BLN55, WL10);
sram_cell_6t_3 inst_cell_9_55 ( BL55, BLN55, WL9);
sram_cell_6t_3 inst_cell_8_55 ( BL55, BLN55, WL8);
sram_cell_6t_3 inst_cell_7_55 ( BL55, BLN55, WL7);
sram_cell_6t_3 inst_cell_6_55 ( BL55, BLN55, WL6);
sram_cell_6t_3 inst_cell_5_55 ( BL55, BLN55, WL5);
sram_cell_6t_3 inst_cell_4_55 ( BL55, BLN55, WL4);
sram_cell_6t_3 inst_cell_3_55 ( BL55, BLN55, WL3);
sram_cell_6t_3 inst_cell_2_55 ( BL55, BLN55, WL2);
sram_cell_6t_3 inst_cell_1_55 ( BL55, BLN55, WL1);
sram_cell_6t_3 inst_cell_0_55 ( BL55, BLN55, WL0);
sram_cell_6t_3 inst_cell_13_54 ( BL54, BLN54, WL13);
sram_cell_6t_3 inst_cell_12_54 ( BL54, BLN54, WL12);
sram_cell_6t_3 inst_cell_11_54 ( BL54, BLN54, WL11);
sram_cell_6t_3 inst_cell_10_54 ( BL54, BLN54, WL10);
sram_cell_6t_3 inst_cell_9_54 ( BL54, BLN54, WL9);
sram_cell_6t_3 inst_cell_8_54 ( BL54, BLN54, WL8);
sram_cell_6t_3 inst_cell_7_54 ( BL54, BLN54, WL7);
sram_cell_6t_3 inst_cell_6_54 ( BL54, BLN54, WL6);
sram_cell_6t_3 inst_cell_5_54 ( BL54, BLN54, WL5);
sram_cell_6t_3 inst_cell_4_54 ( BL54, BLN54, WL4);
sram_cell_6t_3 inst_cell_3_54 ( BL54, BLN54, WL3);
sram_cell_6t_3 inst_cell_2_54 ( BL54, BLN54, WL2);
sram_cell_6t_3 inst_cell_1_54 ( BL54, BLN54, WL1);
sram_cell_6t_3 inst_cell_0_54 ( BL54, BLN54, WL0);
sram_cell_6t_3 inst_cell_13_53 ( BL53, BLN53, WL13);
sram_cell_6t_3 inst_cell_12_53 ( BL53, BLN53, WL12);
sram_cell_6t_3 inst_cell_11_53 ( BL53, BLN53, WL11);
sram_cell_6t_3 inst_cell_10_53 ( BL53, BLN53, WL10);
sram_cell_6t_3 inst_cell_9_53 ( BL53, BLN53, WL9);
sram_cell_6t_3 inst_cell_8_53 ( BL53, BLN53, WL8);
sram_cell_6t_3 inst_cell_7_53 ( BL53, BLN53, WL7);
sram_cell_6t_3 inst_cell_6_53 ( BL53, BLN53, WL6);
sram_cell_6t_3 inst_cell_5_53 ( BL53, BLN53, WL5);
sram_cell_6t_3 inst_cell_4_53 ( BL53, BLN53, WL4);
sram_cell_6t_3 inst_cell_3_53 ( BL53, BLN53, WL3);
sram_cell_6t_3 inst_cell_2_53 ( BL53, BLN53, WL2);
sram_cell_6t_3 inst_cell_1_53 ( BL53, BLN53, WL1);
sram_cell_6t_3 inst_cell_0_53 ( BL53, BLN53, WL0);
sram_cell_6t_3 inst_cell_13_52 ( BL52, BLN52, WL13);
sram_cell_6t_3 inst_cell_12_52 ( BL52, BLN52, WL12);
sram_cell_6t_3 inst_cell_11_52 ( BL52, BLN52, WL11);
sram_cell_6t_3 inst_cell_10_52 ( BL52, BLN52, WL10);
sram_cell_6t_3 inst_cell_9_52 ( BL52, BLN52, WL9);
sram_cell_6t_3 inst_cell_8_52 ( BL52, BLN52, WL8);
sram_cell_6t_3 inst_cell_7_52 ( BL52, BLN52, WL7);
sram_cell_6t_3 inst_cell_6_52 ( BL52, BLN52, WL6);
sram_cell_6t_3 inst_cell_5_52 ( BL52, BLN52, WL5);
sram_cell_6t_3 inst_cell_4_52 ( BL52, BLN52, WL4);
sram_cell_6t_3 inst_cell_3_52 ( BL52, BLN52, WL3);
sram_cell_6t_3 inst_cell_2_52 ( BL52, BLN52, WL2);
sram_cell_6t_3 inst_cell_1_52 ( BL52, BLN52, WL1);
sram_cell_6t_3 inst_cell_0_52 ( BL52, BLN52, WL0);
sram_cell_6t_3 inst_cell_13_51 ( BL51, BLN51, WL13);
sram_cell_6t_3 inst_cell_12_51 ( BL51, BLN51, WL12);
sram_cell_6t_3 inst_cell_11_51 ( BL51, BLN51, WL11);
sram_cell_6t_3 inst_cell_10_51 ( BL51, BLN51, WL10);
sram_cell_6t_3 inst_cell_9_51 ( BL51, BLN51, WL9);
sram_cell_6t_3 inst_cell_8_51 ( BL51, BLN51, WL8);
sram_cell_6t_3 inst_cell_7_51 ( BL51, BLN51, WL7);
sram_cell_6t_3 inst_cell_6_51 ( BL51, BLN51, WL6);
sram_cell_6t_3 inst_cell_5_51 ( BL51, BLN51, WL5);
sram_cell_6t_3 inst_cell_4_51 ( BL51, BLN51, WL4);
sram_cell_6t_3 inst_cell_3_51 ( BL51, BLN51, WL3);
sram_cell_6t_3 inst_cell_2_51 ( BL51, BLN51, WL2);
sram_cell_6t_3 inst_cell_1_51 ( BL51, BLN51, WL1);
sram_cell_6t_3 inst_cell_0_51 ( BL51, BLN51, WL0);
sram_cell_6t_3 inst_cell_13_50 ( BL50, BLN50, WL13);
sram_cell_6t_3 inst_cell_12_50 ( BL50, BLN50, WL12);
sram_cell_6t_3 inst_cell_11_50 ( BL50, BLN50, WL11);
sram_cell_6t_3 inst_cell_10_50 ( BL50, BLN50, WL10);
sram_cell_6t_3 inst_cell_9_50 ( BL50, BLN50, WL9);
sram_cell_6t_3 inst_cell_8_50 ( BL50, BLN50, WL8);
sram_cell_6t_3 inst_cell_7_50 ( BL50, BLN50, WL7);
sram_cell_6t_3 inst_cell_6_50 ( BL50, BLN50, WL6);
sram_cell_6t_3 inst_cell_5_50 ( BL50, BLN50, WL5);
sram_cell_6t_3 inst_cell_4_50 ( BL50, BLN50, WL4);
sram_cell_6t_3 inst_cell_3_50 ( BL50, BLN50, WL3);
sram_cell_6t_3 inst_cell_2_50 ( BL50, BLN50, WL2);
sram_cell_6t_3 inst_cell_1_50 ( BL50, BLN50, WL1);
sram_cell_6t_3 inst_cell_0_50 ( BL50, BLN50, WL0);
sram_cell_6t_3 inst_cell_13_49 ( BL49, BLN49, WL13);
sram_cell_6t_3 inst_cell_12_49 ( BL49, BLN49, WL12);
sram_cell_6t_3 inst_cell_11_49 ( BL49, BLN49, WL11);
sram_cell_6t_3 inst_cell_10_49 ( BL49, BLN49, WL10);
sram_cell_6t_3 inst_cell_9_49 ( BL49, BLN49, WL9);
sram_cell_6t_3 inst_cell_8_49 ( BL49, BLN49, WL8);
sram_cell_6t_3 inst_cell_7_49 ( BL49, BLN49, WL7);
sram_cell_6t_3 inst_cell_6_49 ( BL49, BLN49, WL6);
sram_cell_6t_3 inst_cell_5_49 ( BL49, BLN49, WL5);
sram_cell_6t_3 inst_cell_4_49 ( BL49, BLN49, WL4);
sram_cell_6t_3 inst_cell_3_49 ( BL49, BLN49, WL3);
sram_cell_6t_3 inst_cell_2_49 ( BL49, BLN49, WL2);
sram_cell_6t_3 inst_cell_1_49 ( BL49, BLN49, WL1);
sram_cell_6t_3 inst_cell_0_49 ( BL49, BLN49, WL0);
sram_cell_6t_3 inst_cell_13_48 ( BL48, BLN48, WL13);
sram_cell_6t_3 inst_cell_12_48 ( BL48, BLN48, WL12);
sram_cell_6t_3 inst_cell_11_48 ( BL48, BLN48, WL11);
sram_cell_6t_3 inst_cell_10_48 ( BL48, BLN48, WL10);
sram_cell_6t_3 inst_cell_9_48 ( BL48, BLN48, WL9);
sram_cell_6t_3 inst_cell_8_48 ( BL48, BLN48, WL8);
sram_cell_6t_3 inst_cell_7_48 ( BL48, BLN48, WL7);
sram_cell_6t_3 inst_cell_6_48 ( BL48, BLN48, WL6);
sram_cell_6t_3 inst_cell_5_48 ( BL48, BLN48, WL5);
sram_cell_6t_3 inst_cell_4_48 ( BL48, BLN48, WL4);
sram_cell_6t_3 inst_cell_3_48 ( BL48, BLN48, WL3);
sram_cell_6t_3 inst_cell_2_48 ( BL48, BLN48, WL2);
sram_cell_6t_3 inst_cell_1_48 ( BL48, BLN48, WL1);
sram_cell_6t_3 inst_cell_0_48 ( BL48, BLN48, WL0);
sram_cell_6t_3 inst_cell_13_47 ( BL47, BLN47, WL13);
sram_cell_6t_3 inst_cell_12_47 ( BL47, BLN47, WL12);
sram_cell_6t_3 inst_cell_11_47 ( BL47, BLN47, WL11);
sram_cell_6t_3 inst_cell_10_47 ( BL47, BLN47, WL10);
sram_cell_6t_3 inst_cell_9_47 ( BL47, BLN47, WL9);
sram_cell_6t_3 inst_cell_8_47 ( BL47, BLN47, WL8);
sram_cell_6t_3 inst_cell_7_47 ( BL47, BLN47, WL7);
sram_cell_6t_3 inst_cell_6_47 ( BL47, BLN47, WL6);
sram_cell_6t_3 inst_cell_5_47 ( BL47, BLN47, WL5);
sram_cell_6t_3 inst_cell_4_47 ( BL47, BLN47, WL4);
sram_cell_6t_3 inst_cell_3_47 ( BL47, BLN47, WL3);
sram_cell_6t_3 inst_cell_2_47 ( BL47, BLN47, WL2);
sram_cell_6t_3 inst_cell_1_47 ( BL47, BLN47, WL1);
sram_cell_6t_3 inst_cell_0_47 ( BL47, BLN47, WL0);
sram_cell_6t_3 inst_cell_13_46 ( BL46, BLN46, WL13);
sram_cell_6t_3 inst_cell_12_46 ( BL46, BLN46, WL12);
sram_cell_6t_3 inst_cell_11_46 ( BL46, BLN46, WL11);
sram_cell_6t_3 inst_cell_10_46 ( BL46, BLN46, WL10);
sram_cell_6t_3 inst_cell_9_46 ( BL46, BLN46, WL9);
sram_cell_6t_3 inst_cell_8_46 ( BL46, BLN46, WL8);
sram_cell_6t_3 inst_cell_7_46 ( BL46, BLN46, WL7);
sram_cell_6t_3 inst_cell_6_46 ( BL46, BLN46, WL6);
sram_cell_6t_3 inst_cell_5_46 ( BL46, BLN46, WL5);
sram_cell_6t_3 inst_cell_4_46 ( BL46, BLN46, WL4);
sram_cell_6t_3 inst_cell_3_46 ( BL46, BLN46, WL3);
sram_cell_6t_3 inst_cell_2_46 ( BL46, BLN46, WL2);
sram_cell_6t_3 inst_cell_1_46 ( BL46, BLN46, WL1);
sram_cell_6t_3 inst_cell_0_46 ( BL46, BLN46, WL0);
sram_cell_6t_3 inst_cell_13_45 ( BL45, BLN45, WL13);
sram_cell_6t_3 inst_cell_12_45 ( BL45, BLN45, WL12);
sram_cell_6t_3 inst_cell_11_45 ( BL45, BLN45, WL11);
sram_cell_6t_3 inst_cell_10_45 ( BL45, BLN45, WL10);
sram_cell_6t_3 inst_cell_9_45 ( BL45, BLN45, WL9);
sram_cell_6t_3 inst_cell_8_45 ( BL45, BLN45, WL8);
sram_cell_6t_3 inst_cell_7_45 ( BL45, BLN45, WL7);
sram_cell_6t_3 inst_cell_6_45 ( BL45, BLN45, WL6);
sram_cell_6t_3 inst_cell_5_45 ( BL45, BLN45, WL5);
sram_cell_6t_3 inst_cell_4_45 ( BL45, BLN45, WL4);
sram_cell_6t_3 inst_cell_3_45 ( BL45, BLN45, WL3);
sram_cell_6t_3 inst_cell_2_45 ( BL45, BLN45, WL2);
sram_cell_6t_3 inst_cell_1_45 ( BL45, BLN45, WL1);
sram_cell_6t_3 inst_cell_0_45 ( BL45, BLN45, WL0);
sram_cell_6t_3 inst_cell_13_44 ( BL44, BLN44, WL13);
sram_cell_6t_3 inst_cell_12_44 ( BL44, BLN44, WL12);
sram_cell_6t_3 inst_cell_11_44 ( BL44, BLN44, WL11);
sram_cell_6t_3 inst_cell_10_44 ( BL44, BLN44, WL10);
sram_cell_6t_3 inst_cell_9_44 ( BL44, BLN44, WL9);
sram_cell_6t_3 inst_cell_8_44 ( BL44, BLN44, WL8);
sram_cell_6t_3 inst_cell_7_44 ( BL44, BLN44, WL7);
sram_cell_6t_3 inst_cell_6_44 ( BL44, BLN44, WL6);
sram_cell_6t_3 inst_cell_5_44 ( BL44, BLN44, WL5);
sram_cell_6t_3 inst_cell_4_44 ( BL44, BLN44, WL4);
sram_cell_6t_3 inst_cell_3_44 ( BL44, BLN44, WL3);
sram_cell_6t_3 inst_cell_2_44 ( BL44, BLN44, WL2);
sram_cell_6t_3 inst_cell_1_44 ( BL44, BLN44, WL1);
sram_cell_6t_3 inst_cell_0_44 ( BL44, BLN44, WL0);
sram_cell_6t_3 inst_cell_13_43 ( BL43, BLN43, WL13);
sram_cell_6t_3 inst_cell_12_43 ( BL43, BLN43, WL12);
sram_cell_6t_3 inst_cell_11_43 ( BL43, BLN43, WL11);
sram_cell_6t_3 inst_cell_10_43 ( BL43, BLN43, WL10);
sram_cell_6t_3 inst_cell_9_43 ( BL43, BLN43, WL9);
sram_cell_6t_3 inst_cell_8_43 ( BL43, BLN43, WL8);
sram_cell_6t_3 inst_cell_7_43 ( BL43, BLN43, WL7);
sram_cell_6t_3 inst_cell_6_43 ( BL43, BLN43, WL6);
sram_cell_6t_3 inst_cell_5_43 ( BL43, BLN43, WL5);
sram_cell_6t_3 inst_cell_4_43 ( BL43, BLN43, WL4);
sram_cell_6t_3 inst_cell_3_43 ( BL43, BLN43, WL3);
sram_cell_6t_3 inst_cell_2_43 ( BL43, BLN43, WL2);
sram_cell_6t_3 inst_cell_1_43 ( BL43, BLN43, WL1);
sram_cell_6t_3 inst_cell_0_43 ( BL43, BLN43, WL0);
sram_cell_6t_3 inst_cell_13_42 ( BL42, BLN42, WL13);
sram_cell_6t_3 inst_cell_12_42 ( BL42, BLN42, WL12);
sram_cell_6t_3 inst_cell_11_42 ( BL42, BLN42, WL11);
sram_cell_6t_3 inst_cell_10_42 ( BL42, BLN42, WL10);
sram_cell_6t_3 inst_cell_9_42 ( BL42, BLN42, WL9);
sram_cell_6t_3 inst_cell_8_42 ( BL42, BLN42, WL8);
sram_cell_6t_3 inst_cell_7_42 ( BL42, BLN42, WL7);
sram_cell_6t_3 inst_cell_6_42 ( BL42, BLN42, WL6);
sram_cell_6t_3 inst_cell_5_42 ( BL42, BLN42, WL5);
sram_cell_6t_3 inst_cell_4_42 ( BL42, BLN42, WL4);
sram_cell_6t_3 inst_cell_3_42 ( BL42, BLN42, WL3);
sram_cell_6t_3 inst_cell_2_42 ( BL42, BLN42, WL2);
sram_cell_6t_3 inst_cell_1_42 ( BL42, BLN42, WL1);
sram_cell_6t_3 inst_cell_0_42 ( BL42, BLN42, WL0);
sram_cell_6t_3 inst_cell_13_41 ( BL41, BLN41, WL13);
sram_cell_6t_3 inst_cell_12_41 ( BL41, BLN41, WL12);
sram_cell_6t_3 inst_cell_11_41 ( BL41, BLN41, WL11);
sram_cell_6t_3 inst_cell_10_41 ( BL41, BLN41, WL10);
sram_cell_6t_3 inst_cell_9_41 ( BL41, BLN41, WL9);
sram_cell_6t_3 inst_cell_8_41 ( BL41, BLN41, WL8);
sram_cell_6t_3 inst_cell_7_41 ( BL41, BLN41, WL7);
sram_cell_6t_3 inst_cell_6_41 ( BL41, BLN41, WL6);
sram_cell_6t_3 inst_cell_5_41 ( BL41, BLN41, WL5);
sram_cell_6t_3 inst_cell_4_41 ( BL41, BLN41, WL4);
sram_cell_6t_3 inst_cell_3_41 ( BL41, BLN41, WL3);
sram_cell_6t_3 inst_cell_2_41 ( BL41, BLN41, WL2);
sram_cell_6t_3 inst_cell_1_41 ( BL41, BLN41, WL1);
sram_cell_6t_3 inst_cell_0_41 ( BL41, BLN41, WL0);
sram_cell_6t_3 inst_cell_13_40 ( BL40, BLN40, WL13);
sram_cell_6t_3 inst_cell_12_40 ( BL40, BLN40, WL12);
sram_cell_6t_3 inst_cell_11_40 ( BL40, BLN40, WL11);
sram_cell_6t_3 inst_cell_10_40 ( BL40, BLN40, WL10);
sram_cell_6t_3 inst_cell_9_40 ( BL40, BLN40, WL9);
sram_cell_6t_3 inst_cell_8_40 ( BL40, BLN40, WL8);
sram_cell_6t_3 inst_cell_7_40 ( BL40, BLN40, WL7);
sram_cell_6t_3 inst_cell_6_40 ( BL40, BLN40, WL6);
sram_cell_6t_3 inst_cell_5_40 ( BL40, BLN40, WL5);
sram_cell_6t_3 inst_cell_4_40 ( BL40, BLN40, WL4);
sram_cell_6t_3 inst_cell_3_40 ( BL40, BLN40, WL3);
sram_cell_6t_3 inst_cell_2_40 ( BL40, BLN40, WL2);
sram_cell_6t_3 inst_cell_1_40 ( BL40, BLN40, WL1);
sram_cell_6t_3 inst_cell_0_40 ( BL40, BLN40, WL0);
sram_cell_6t_3 inst_cell_13_39 ( BL39, BLN39, WL13);
sram_cell_6t_3 inst_cell_12_39 ( BL39, BLN39, WL12);
sram_cell_6t_3 inst_cell_11_39 ( BL39, BLN39, WL11);
sram_cell_6t_3 inst_cell_10_39 ( BL39, BLN39, WL10);
sram_cell_6t_3 inst_cell_9_39 ( BL39, BLN39, WL9);
sram_cell_6t_3 inst_cell_8_39 ( BL39, BLN39, WL8);
sram_cell_6t_3 inst_cell_7_39 ( BL39, BLN39, WL7);
sram_cell_6t_3 inst_cell_6_39 ( BL39, BLN39, WL6);
sram_cell_6t_3 inst_cell_5_39 ( BL39, BLN39, WL5);
sram_cell_6t_3 inst_cell_4_39 ( BL39, BLN39, WL4);
sram_cell_6t_3 inst_cell_3_39 ( BL39, BLN39, WL3);
sram_cell_6t_3 inst_cell_2_39 ( BL39, BLN39, WL2);
sram_cell_6t_3 inst_cell_1_39 ( BL39, BLN39, WL1);
sram_cell_6t_3 inst_cell_0_39 ( BL39, BLN39, WL0);
sram_cell_6t_3 inst_cell_13_38 ( BL38, BLN38, WL13);
sram_cell_6t_3 inst_cell_12_38 ( BL38, BLN38, WL12);
sram_cell_6t_3 inst_cell_11_38 ( BL38, BLN38, WL11);
sram_cell_6t_3 inst_cell_10_38 ( BL38, BLN38, WL10);
sram_cell_6t_3 inst_cell_9_38 ( BL38, BLN38, WL9);
sram_cell_6t_3 inst_cell_8_38 ( BL38, BLN38, WL8);
sram_cell_6t_3 inst_cell_7_38 ( BL38, BLN38, WL7);
sram_cell_6t_3 inst_cell_6_38 ( BL38, BLN38, WL6);
sram_cell_6t_3 inst_cell_5_38 ( BL38, BLN38, WL5);
sram_cell_6t_3 inst_cell_4_38 ( BL38, BLN38, WL4);
sram_cell_6t_3 inst_cell_3_38 ( BL38, BLN38, WL3);
sram_cell_6t_3 inst_cell_2_38 ( BL38, BLN38, WL2);
sram_cell_6t_3 inst_cell_1_38 ( BL38, BLN38, WL1);
sram_cell_6t_3 inst_cell_0_38 ( BL38, BLN38, WL0);
sram_cell_6t_3 inst_cell_13_37 ( BL37, BLN37, WL13);
sram_cell_6t_3 inst_cell_12_37 ( BL37, BLN37, WL12);
sram_cell_6t_3 inst_cell_11_37 ( BL37, BLN37, WL11);
sram_cell_6t_3 inst_cell_10_37 ( BL37, BLN37, WL10);
sram_cell_6t_3 inst_cell_9_37 ( BL37, BLN37, WL9);
sram_cell_6t_3 inst_cell_8_37 ( BL37, BLN37, WL8);
sram_cell_6t_3 inst_cell_7_37 ( BL37, BLN37, WL7);
sram_cell_6t_3 inst_cell_6_37 ( BL37, BLN37, WL6);
sram_cell_6t_3 inst_cell_5_37 ( BL37, BLN37, WL5);
sram_cell_6t_3 inst_cell_4_37 ( BL37, BLN37, WL4);
sram_cell_6t_3 inst_cell_3_37 ( BL37, BLN37, WL3);
sram_cell_6t_3 inst_cell_2_37 ( BL37, BLN37, WL2);
sram_cell_6t_3 inst_cell_1_37 ( BL37, BLN37, WL1);
sram_cell_6t_3 inst_cell_0_37 ( BL37, BLN37, WL0);
sram_cell_6t_3 inst_cell_13_36 ( BL36, BLN36, WL13);
sram_cell_6t_3 inst_cell_12_36 ( BL36, BLN36, WL12);
sram_cell_6t_3 inst_cell_11_36 ( BL36, BLN36, WL11);
sram_cell_6t_3 inst_cell_10_36 ( BL36, BLN36, WL10);
sram_cell_6t_3 inst_cell_9_36 ( BL36, BLN36, WL9);
sram_cell_6t_3 inst_cell_8_36 ( BL36, BLN36, WL8);
sram_cell_6t_3 inst_cell_7_36 ( BL36, BLN36, WL7);
sram_cell_6t_3 inst_cell_6_36 ( BL36, BLN36, WL6);
sram_cell_6t_3 inst_cell_5_36 ( BL36, BLN36, WL5);
sram_cell_6t_3 inst_cell_4_36 ( BL36, BLN36, WL4);
sram_cell_6t_3 inst_cell_3_36 ( BL36, BLN36, WL3);
sram_cell_6t_3 inst_cell_2_36 ( BL36, BLN36, WL2);
sram_cell_6t_3 inst_cell_1_36 ( BL36, BLN36, WL1);
sram_cell_6t_3 inst_cell_0_36 ( BL36, BLN36, WL0);
sram_cell_6t_3 inst_cell_13_35 ( BL35, BLN35, WL13);
sram_cell_6t_3 inst_cell_12_35 ( BL35, BLN35, WL12);
sram_cell_6t_3 inst_cell_11_35 ( BL35, BLN35, WL11);
sram_cell_6t_3 inst_cell_10_35 ( BL35, BLN35, WL10);
sram_cell_6t_3 inst_cell_9_35 ( BL35, BLN35, WL9);
sram_cell_6t_3 inst_cell_8_35 ( BL35, BLN35, WL8);
sram_cell_6t_3 inst_cell_7_35 ( BL35, BLN35, WL7);
sram_cell_6t_3 inst_cell_6_35 ( BL35, BLN35, WL6);
sram_cell_6t_3 inst_cell_5_35 ( BL35, BLN35, WL5);
sram_cell_6t_3 inst_cell_4_35 ( BL35, BLN35, WL4);
sram_cell_6t_3 inst_cell_3_35 ( BL35, BLN35, WL3);
sram_cell_6t_3 inst_cell_2_35 ( BL35, BLN35, WL2);
sram_cell_6t_3 inst_cell_1_35 ( BL35, BLN35, WL1);
sram_cell_6t_3 inst_cell_0_35 ( BL35, BLN35, WL0);
sram_cell_6t_3 inst_cell_13_34 ( BL34, BLN34, WL13);
sram_cell_6t_3 inst_cell_12_34 ( BL34, BLN34, WL12);
sram_cell_6t_3 inst_cell_11_34 ( BL34, BLN34, WL11);
sram_cell_6t_3 inst_cell_10_34 ( BL34, BLN34, WL10);
sram_cell_6t_3 inst_cell_9_34 ( BL34, BLN34, WL9);
sram_cell_6t_3 inst_cell_8_34 ( BL34, BLN34, WL8);
sram_cell_6t_3 inst_cell_7_34 ( BL34, BLN34, WL7);
sram_cell_6t_3 inst_cell_6_34 ( BL34, BLN34, WL6);
sram_cell_6t_3 inst_cell_5_34 ( BL34, BLN34, WL5);
sram_cell_6t_3 inst_cell_4_34 ( BL34, BLN34, WL4);
sram_cell_6t_3 inst_cell_3_34 ( BL34, BLN34, WL3);
sram_cell_6t_3 inst_cell_2_34 ( BL34, BLN34, WL2);
sram_cell_6t_3 inst_cell_1_34 ( BL34, BLN34, WL1);
sram_cell_6t_3 inst_cell_0_34 ( BL34, BLN34, WL0);
sram_cell_6t_3 inst_cell_13_33 ( BL33, BLN33, WL13);
sram_cell_6t_3 inst_cell_12_33 ( BL33, BLN33, WL12);
sram_cell_6t_3 inst_cell_11_33 ( BL33, BLN33, WL11);
sram_cell_6t_3 inst_cell_10_33 ( BL33, BLN33, WL10);
sram_cell_6t_3 inst_cell_9_33 ( BL33, BLN33, WL9);
sram_cell_6t_3 inst_cell_8_33 ( BL33, BLN33, WL8);
sram_cell_6t_3 inst_cell_7_33 ( BL33, BLN33, WL7);
sram_cell_6t_3 inst_cell_6_33 ( BL33, BLN33, WL6);
sram_cell_6t_3 inst_cell_5_33 ( BL33, BLN33, WL5);
sram_cell_6t_3 inst_cell_4_33 ( BL33, BLN33, WL4);
sram_cell_6t_3 inst_cell_3_33 ( BL33, BLN33, WL3);
sram_cell_6t_3 inst_cell_2_33 ( BL33, BLN33, WL2);
sram_cell_6t_3 inst_cell_1_33 ( BL33, BLN33, WL1);
sram_cell_6t_3 inst_cell_0_33 ( BL33, BLN33, WL0);
sram_cell_6t_3 inst_cell_13_32 ( BL32, BLN32, WL13);
sram_cell_6t_3 inst_cell_12_32 ( BL32, BLN32, WL12);
sram_cell_6t_3 inst_cell_11_32 ( BL32, BLN32, WL11);
sram_cell_6t_3 inst_cell_10_32 ( BL32, BLN32, WL10);
sram_cell_6t_3 inst_cell_9_32 ( BL32, BLN32, WL9);
sram_cell_6t_3 inst_cell_8_32 ( BL32, BLN32, WL8);
sram_cell_6t_3 inst_cell_7_32 ( BL32, BLN32, WL7);
sram_cell_6t_3 inst_cell_6_32 ( BL32, BLN32, WL6);
sram_cell_6t_3 inst_cell_5_32 ( BL32, BLN32, WL5);
sram_cell_6t_3 inst_cell_4_32 ( BL32, BLN32, WL4);
sram_cell_6t_3 inst_cell_3_32 ( BL32, BLN32, WL3);
sram_cell_6t_3 inst_cell_2_32 ( BL32, BLN32, WL2);
sram_cell_6t_3 inst_cell_1_32 ( BL32, BLN32, WL1);
sram_cell_6t_3 inst_cell_0_32 ( BL32, BLN32, WL0);
sram_cell_6t_3 inst_cell_13_31 ( BL31, BLN31, WL13);
sram_cell_6t_3 inst_cell_12_31 ( BL31, BLN31, WL12);
sram_cell_6t_3 inst_cell_11_31 ( BL31, BLN31, WL11);
sram_cell_6t_3 inst_cell_10_31 ( BL31, BLN31, WL10);
sram_cell_6t_3 inst_cell_9_31 ( BL31, BLN31, WL9);
sram_cell_6t_3 inst_cell_8_31 ( BL31, BLN31, WL8);
sram_cell_6t_3 inst_cell_7_31 ( BL31, BLN31, WL7);
sram_cell_6t_3 inst_cell_6_31 ( BL31, BLN31, WL6);
sram_cell_6t_3 inst_cell_5_31 ( BL31, BLN31, WL5);
sram_cell_6t_3 inst_cell_4_31 ( BL31, BLN31, WL4);
sram_cell_6t_3 inst_cell_3_31 ( BL31, BLN31, WL3);
sram_cell_6t_3 inst_cell_2_31 ( BL31, BLN31, WL2);
sram_cell_6t_3 inst_cell_1_31 ( BL31, BLN31, WL1);
sram_cell_6t_3 inst_cell_0_31 ( BL31, BLN31, WL0);
sram_cell_6t_3 inst_cell_13_30 ( BL30, BLN30, WL13);
sram_cell_6t_3 inst_cell_12_30 ( BL30, BLN30, WL12);
sram_cell_6t_3 inst_cell_11_30 ( BL30, BLN30, WL11);
sram_cell_6t_3 inst_cell_10_30 ( BL30, BLN30, WL10);
sram_cell_6t_3 inst_cell_9_30 ( BL30, BLN30, WL9);
sram_cell_6t_3 inst_cell_8_30 ( BL30, BLN30, WL8);
sram_cell_6t_3 inst_cell_7_30 ( BL30, BLN30, WL7);
sram_cell_6t_3 inst_cell_6_30 ( BL30, BLN30, WL6);
sram_cell_6t_3 inst_cell_5_30 ( BL30, BLN30, WL5);
sram_cell_6t_3 inst_cell_4_30 ( BL30, BLN30, WL4);
sram_cell_6t_3 inst_cell_3_30 ( BL30, BLN30, WL3);
sram_cell_6t_3 inst_cell_2_30 ( BL30, BLN30, WL2);
sram_cell_6t_3 inst_cell_1_30 ( BL30, BLN30, WL1);
sram_cell_6t_3 inst_cell_0_30 ( BL30, BLN30, WL0);
sram_cell_6t_3 inst_cell_13_29 ( BL29, BLN29, WL13);
sram_cell_6t_3 inst_cell_12_29 ( BL29, BLN29, WL12);
sram_cell_6t_3 inst_cell_11_29 ( BL29, BLN29, WL11);
sram_cell_6t_3 inst_cell_10_29 ( BL29, BLN29, WL10);
sram_cell_6t_3 inst_cell_9_29 ( BL29, BLN29, WL9);
sram_cell_6t_3 inst_cell_8_29 ( BL29, BLN29, WL8);
sram_cell_6t_3 inst_cell_7_29 ( BL29, BLN29, WL7);
sram_cell_6t_3 inst_cell_6_29 ( BL29, BLN29, WL6);
sram_cell_6t_3 inst_cell_13_28 ( BL28, BLN28, WL13);
sram_cell_6t_3 inst_cell_12_28 ( BL28, BLN28, WL12);
sram_cell_6t_3 inst_cell_11_28 ( BL28, BLN28, WL11);
sram_cell_6t_3 inst_cell_10_28 ( BL28, BLN28, WL10);
sram_cell_6t_3 inst_cell_9_28 ( BL28, BLN28, WL9);
sram_cell_6t_3 inst_cell_8_28 ( BL28, BLN28, WL8);
sram_cell_6t_3 inst_cell_7_28 ( BL28, BLN28, WL7);
sram_cell_6t_3 inst_cell_6_28 ( BL28, BLN28, WL6);
sram_cell_6t_3 inst_cell_5_28 ( BL28, BLN28, WL5);
sram_cell_6t_3 inst_cell_4_28 ( BL28, BLN28, WL4);
sram_cell_6t_3 inst_cell_3_28 ( BL28, BLN28, WL3);
sram_cell_6t_3 inst_cell_2_28 ( BL28, BLN28, WL2);
sram_cell_6t_3 inst_cell_1_28 ( BL28, BLN28, WL1);
sram_cell_6t_3 inst_cell_0_28 ( BL28, BLN28, WL0);
sram_cell_6t_3 inst_cell_13_27 ( BL27, BLN27, WL13);
sram_cell_6t_3 inst_cell_12_27 ( BL27, BLN27, WL12);
sram_cell_6t_3 inst_cell_11_27 ( BL27, BLN27, WL11);
sram_cell_6t_3 inst_cell_10_27 ( BL27, BLN27, WL10);
sram_cell_6t_3 inst_cell_9_27 ( BL27, BLN27, WL9);
sram_cell_6t_3 inst_cell_8_27 ( BL27, BLN27, WL8);
sram_cell_6t_3 inst_cell_7_27 ( BL27, BLN27, WL7);
sram_cell_6t_3 inst_cell_6_27 ( BL27, BLN27, WL6);
sram_cell_6t_3 inst_cell_5_27 ( BL27, BLN27, WL5);
sram_cell_6t_3 inst_cell_4_27 ( BL27, BLN27, WL4);
sram_cell_6t_3 inst_cell_3_27 ( BL27, BLN27, WL3);
sram_cell_6t_3 inst_cell_2_27 ( BL27, BLN27, WL2);
sram_cell_6t_3 inst_cell_1_27 ( BL27, BLN27, WL1);
sram_cell_6t_3 inst_cell_0_27 ( BL27, BLN27, WL0);
sram_cell_6t_3 inst_cell_13_26 ( BL26, BLN26, WL13);
sram_cell_6t_3 inst_cell_12_26 ( BL26, BLN26, WL12);
sram_cell_6t_3 inst_cell_11_26 ( BL26, BLN26, WL11);
sram_cell_6t_3 inst_cell_10_26 ( BL26, BLN26, WL10);
sram_cell_6t_3 inst_cell_9_26 ( BL26, BLN26, WL9);
sram_cell_6t_3 inst_cell_8_26 ( BL26, BLN26, WL8);
sram_cell_6t_3 inst_cell_7_26 ( BL26, BLN26, WL7);
sram_cell_6t_3 inst_cell_6_26 ( BL26, BLN26, WL6);
sram_cell_6t_3 inst_cell_5_26 ( BL26, BLN26, WL5);
sram_cell_6t_3 inst_cell_4_26 ( BL26, BLN26, WL4);
sram_cell_6t_3 inst_cell_3_26 ( BL26, BLN26, WL3);
sram_cell_6t_3 inst_cell_2_26 ( BL26, BLN26, WL2);
sram_cell_6t_3 inst_cell_1_26 ( BL26, BLN26, WL1);
sram_cell_6t_3 inst_cell_0_26 ( BL26, BLN26, WL0);
sram_cell_6t_3 inst_cell_13_25 ( BL25, BLN25, WL13);
sram_cell_6t_3 inst_cell_12_25 ( BL25, BLN25, WL12);
sram_cell_6t_3 inst_cell_11_25 ( BL25, BLN25, WL11);
sram_cell_6t_3 inst_cell_10_25 ( BL25, BLN25, WL10);
sram_cell_6t_3 inst_cell_9_25 ( BL25, BLN25, WL9);
sram_cell_6t_3 inst_cell_8_25 ( BL25, BLN25, WL8);
sram_cell_6t_3 inst_cell_7_25 ( BL25, BLN25, WL7);
sram_cell_6t_3 inst_cell_6_25 ( BL25, BLN25, WL6);
sram_cell_6t_3 inst_cell_5_25 ( BL25, BLN25, WL5);
sram_cell_6t_3 inst_cell_4_25 ( BL25, BLN25, WL4);
sram_cell_6t_3 inst_cell_3_25 ( BL25, BLN25, WL3);
sram_cell_6t_3 inst_cell_2_25 ( BL25, BLN25, WL2);
sram_cell_6t_3 inst_cell_1_25 ( BL25, BLN25, WL1);
sram_cell_6t_3 inst_cell_0_25 ( BL25, BLN25, WL0);
sram_cell_6t_3 inst_cell_13_24 ( BL24, BLN24, WL13);
sram_cell_6t_3 inst_cell_12_24 ( BL24, BLN24, WL12);
sram_cell_6t_3 inst_cell_11_24 ( BL24, BLN24, WL11);
sram_cell_6t_3 inst_cell_10_24 ( BL24, BLN24, WL10);
sram_cell_6t_3 inst_cell_9_24 ( BL24, BLN24, WL9);
sram_cell_6t_3 inst_cell_8_24 ( BL24, BLN24, WL8);
sram_cell_6t_3 inst_cell_7_24 ( BL24, BLN24, WL7);
sram_cell_6t_3 inst_cell_6_24 ( BL24, BLN24, WL6);
sram_cell_6t_3 inst_cell_5_24 ( BL24, BLN24, WL5);
sram_cell_6t_3 inst_cell_4_24 ( BL24, BLN24, WL4);
sram_cell_6t_3 inst_cell_3_24 ( BL24, BLN24, WL3);
sram_cell_6t_3 inst_cell_2_24 ( BL24, BLN24, WL2);
sram_cell_6t_3 inst_cell_1_24 ( BL24, BLN24, WL1);
sram_cell_6t_3 inst_cell_0_24 ( BL24, BLN24, WL0);
sram_cell_6t_3 inst_cell_13_23 ( BL23, BLN23, WL13);
sram_cell_6t_3 inst_cell_12_23 ( BL23, BLN23, WL12);
sram_cell_6t_3 inst_cell_11_23 ( BL23, BLN23, WL11);
sram_cell_6t_3 inst_cell_10_23 ( BL23, BLN23, WL10);
sram_cell_6t_3 inst_cell_9_23 ( BL23, BLN23, WL9);
sram_cell_6t_3 inst_cell_8_23 ( BL23, BLN23, WL8);
sram_cell_6t_3 inst_cell_7_23 ( BL23, BLN23, WL7);
sram_cell_6t_3 inst_cell_6_23 ( BL23, BLN23, WL6);
sram_cell_6t_3 inst_cell_5_23 ( BL23, BLN23, WL5);
sram_cell_6t_3 inst_cell_4_23 ( BL23, BLN23, WL4);
sram_cell_6t_3 inst_cell_3_23 ( BL23, BLN23, WL3);
sram_cell_6t_3 inst_cell_2_23 ( BL23, BLN23, WL2);
sram_cell_6t_3 inst_cell_1_23 ( BL23, BLN23, WL1);
sram_cell_6t_3 inst_cell_0_23 ( BL23, BLN23, WL0);
sram_cell_6t_3 inst_cell_13_22 ( BL22, BLN22, WL13);
sram_cell_6t_3 inst_cell_12_22 ( BL22, BLN22, WL12);
sram_cell_6t_3 inst_cell_11_22 ( BL22, BLN22, WL11);
sram_cell_6t_3 inst_cell_10_22 ( BL22, BLN22, WL10);
sram_cell_6t_3 inst_cell_9_22 ( BL22, BLN22, WL9);
sram_cell_6t_3 inst_cell_8_22 ( BL22, BLN22, WL8);
sram_cell_6t_3 inst_cell_7_22 ( BL22, BLN22, WL7);
sram_cell_6t_3 inst_cell_6_22 ( BL22, BLN22, WL6);
sram_cell_6t_3 inst_cell_5_22 ( BL22, BLN22, WL5);
sram_cell_6t_3 inst_cell_4_22 ( BL22, BLN22, WL4);
sram_cell_6t_3 inst_cell_3_22 ( BL22, BLN22, WL3);
sram_cell_6t_3 inst_cell_2_22 ( BL22, BLN22, WL2);
sram_cell_6t_3 inst_cell_1_22 ( BL22, BLN22, WL1);
sram_cell_6t_3 inst_cell_0_22 ( BL22, BLN22, WL0);
sram_cell_6t_3 inst_cell_13_21 ( BL21, BLN21, WL13);
sram_cell_6t_3 inst_cell_12_21 ( BL21, BLN21, WL12);
sram_cell_6t_3 inst_cell_11_21 ( BL21, BLN21, WL11);
sram_cell_6t_3 inst_cell_10_21 ( BL21, BLN21, WL10);
sram_cell_6t_3 inst_cell_9_21 ( BL21, BLN21, WL9);
sram_cell_6t_3 inst_cell_8_21 ( BL21, BLN21, WL8);
sram_cell_6t_3 inst_cell_7_21 ( BL21, BLN21, WL7);
sram_cell_6t_3 inst_cell_6_21 ( BL21, BLN21, WL6);
sram_cell_6t_3 inst_cell_5_21 ( BL21, BLN21, WL5);
sram_cell_6t_3 inst_cell_4_21 ( BL21, BLN21, WL4);
sram_cell_6t_3 inst_cell_3_21 ( BL21, BLN21, WL3);
sram_cell_6t_3 inst_cell_2_21 ( BL21, BLN21, WL2);
sram_cell_6t_3 inst_cell_1_21 ( BL21, BLN21, WL1);
sram_cell_6t_3 inst_cell_0_21 ( BL21, BLN21, WL0);
sram_cell_6t_3 inst_cell_13_20 ( BL20, BLN20, WL13);
sram_cell_6t_3 inst_cell_12_20 ( BL20, BLN20, WL12);
sram_cell_6t_3 inst_cell_11_20 ( BL20, BLN20, WL11);
sram_cell_6t_3 inst_cell_10_20 ( BL20, BLN20, WL10);
sram_cell_6t_3 inst_cell_9_20 ( BL20, BLN20, WL9);
sram_cell_6t_3 inst_cell_8_20 ( BL20, BLN20, WL8);
sram_cell_6t_3 inst_cell_7_20 ( BL20, BLN20, WL7);
sram_cell_6t_3 inst_cell_6_20 ( BL20, BLN20, WL6);
sram_cell_6t_3 inst_cell_5_20 ( BL20, BLN20, WL5);
sram_cell_6t_3 inst_cell_4_20 ( BL20, BLN20, WL4);
sram_cell_6t_3 inst_cell_3_20 ( BL20, BLN20, WL3);
sram_cell_6t_3 inst_cell_2_20 ( BL20, BLN20, WL2);
sram_cell_6t_3 inst_cell_1_20 ( BL20, BLN20, WL1);
sram_cell_6t_3 inst_cell_0_20 ( BL20, BLN20, WL0);
sram_cell_6t_3 inst_cell_13_19 ( BL19, BLN19, WL13);
sram_cell_6t_3 inst_cell_12_19 ( BL19, BLN19, WL12);
sram_cell_6t_3 inst_cell_11_19 ( BL19, BLN19, WL11);
sram_cell_6t_3 inst_cell_10_19 ( BL19, BLN19, WL10);
sram_cell_6t_3 inst_cell_9_19 ( BL19, BLN19, WL9);
sram_cell_6t_3 inst_cell_8_19 ( BL19, BLN19, WL8);
sram_cell_6t_3 inst_cell_7_19 ( BL19, BLN19, WL7);
sram_cell_6t_3 inst_cell_6_19 ( BL19, BLN19, WL6);
sram_cell_6t_3 inst_cell_5_19 ( BL19, BLN19, WL5);
sram_cell_6t_3 inst_cell_4_19 ( BL19, BLN19, WL4);
sram_cell_6t_3 inst_cell_3_19 ( BL19, BLN19, WL3);
sram_cell_6t_3 inst_cell_2_19 ( BL19, BLN19, WL2);
sram_cell_6t_3 inst_cell_1_19 ( BL19, BLN19, WL1);
sram_cell_6t_3 inst_cell_0_19 ( BL19, BLN19, WL0);
sram_cell_6t_3 inst_cell_13_18 ( BL18, BLN18, WL13);
sram_cell_6t_3 inst_cell_12_18 ( BL18, BLN18, WL12);
sram_cell_6t_3 inst_cell_11_18 ( BL18, BLN18, WL11);
sram_cell_6t_3 inst_cell_10_18 ( BL18, BLN18, WL10);
sram_cell_6t_3 inst_cell_9_18 ( BL18, BLN18, WL9);
sram_cell_6t_3 inst_cell_8_18 ( BL18, BLN18, WL8);
sram_cell_6t_3 inst_cell_7_18 ( BL18, BLN18, WL7);
sram_cell_6t_3 inst_cell_6_18 ( BL18, BLN18, WL6);
sram_cell_6t_3 inst_cell_5_18 ( BL18, BLN18, WL5);
sram_cell_6t_3 inst_cell_4_18 ( BL18, BLN18, WL4);
sram_cell_6t_3 inst_cell_3_18 ( BL18, BLN18, WL3);
sram_cell_6t_3 inst_cell_2_18 ( BL18, BLN18, WL2);
sram_cell_6t_3 inst_cell_1_18 ( BL18, BLN18, WL1);
sram_cell_6t_3 inst_cell_0_18 ( BL18, BLN18, WL0);
sram_cell_6t_3 inst_cell_13_17 ( BL17, BLN17, WL13);
sram_cell_6t_3 inst_cell_12_17 ( BL17, BLN17, WL12);
sram_cell_6t_3 inst_cell_11_17 ( BL17, BLN17, WL11);
sram_cell_6t_3 inst_cell_10_17 ( BL17, BLN17, WL10);
sram_cell_6t_3 inst_cell_9_17 ( BL17, BLN17, WL9);
sram_cell_6t_3 inst_cell_8_17 ( BL17, BLN17, WL8);
sram_cell_6t_3 inst_cell_7_17 ( BL17, BLN17, WL7);
sram_cell_6t_3 inst_cell_6_17 ( BL17, BLN17, WL6);
sram_cell_6t_3 inst_cell_5_17 ( BL17, BLN17, WL5);
sram_cell_6t_3 inst_cell_4_17 ( BL17, BLN17, WL4);
sram_cell_6t_3 inst_cell_3_17 ( BL17, BLN17, WL3);
sram_cell_6t_3 inst_cell_2_17 ( BL17, BLN17, WL2);
sram_cell_6t_3 inst_cell_1_17 ( BL17, BLN17, WL1);
sram_cell_6t_3 inst_cell_0_17 ( BL17, BLN17, WL0);
sram_cell_6t_3 inst_cell_13_16 ( BL16, BLN16, WL13);
sram_cell_6t_3 inst_cell_12_16 ( BL16, BLN16, WL12);
sram_cell_6t_3 inst_cell_11_16 ( BL16, BLN16, WL11);
sram_cell_6t_3 inst_cell_10_16 ( BL16, BLN16, WL10);
sram_cell_6t_3 inst_cell_9_16 ( BL16, BLN16, WL9);
sram_cell_6t_3 inst_cell_8_16 ( BL16, BLN16, WL8);
sram_cell_6t_3 inst_cell_7_16 ( BL16, BLN16, WL7);
sram_cell_6t_3 inst_cell_6_16 ( BL16, BLN16, WL6);
sram_cell_6t_3 inst_cell_5_16 ( BL16, BLN16, WL5);
sram_cell_6t_3 inst_cell_4_16 ( BL16, BLN16, WL4);
sram_cell_6t_3 inst_cell_3_16 ( BL16, BLN16, WL3);
sram_cell_6t_3 inst_cell_2_16 ( BL16, BLN16, WL2);
sram_cell_6t_3 inst_cell_1_16 ( BL16, BLN16, WL1);
sram_cell_6t_3 inst_cell_0_16 ( BL16, BLN16, WL0);
sram_cell_6t_3 inst_cell_13_15 ( BL15, BLN15, WL13);
sram_cell_6t_3 inst_cell_12_15 ( BL15, BLN15, WL12);
sram_cell_6t_3 inst_cell_11_15 ( BL15, BLN15, WL11);
sram_cell_6t_3 inst_cell_10_15 ( BL15, BLN15, WL10);
sram_cell_6t_3 inst_cell_9_15 ( BL15, BLN15, WL9);
sram_cell_6t_3 inst_cell_8_15 ( BL15, BLN15, WL8);
sram_cell_6t_3 inst_cell_7_15 ( BL15, BLN15, WL7);
sram_cell_6t_3 inst_cell_6_15 ( BL15, BLN15, WL6);
sram_cell_6t_3 inst_cell_5_15 ( BL15, BLN15, WL5);
sram_cell_6t_3 inst_cell_4_15 ( BL15, BLN15, WL4);
sram_cell_6t_3 inst_cell_3_15 ( BL15, BLN15, WL3);
sram_cell_6t_3 inst_cell_2_15 ( BL15, BLN15, WL2);
sram_cell_6t_3 inst_cell_1_15 ( BL15, BLN15, WL1);
sram_cell_6t_3 inst_cell_0_15 ( BL15, BLN15, WL0);
sram_cell_6t_3 inst_cell_13_14 ( BL14, BLN14, WL13);
sram_cell_6t_3 inst_cell_12_14 ( BL14, BLN14, WL12);
sram_cell_6t_3 inst_cell_11_14 ( BL14, BLN14, WL11);
sram_cell_6t_3 inst_cell_10_14 ( BL14, BLN14, WL10);
sram_cell_6t_3 inst_cell_9_14 ( BL14, BLN14, WL9);
sram_cell_6t_3 inst_cell_8_14 ( BL14, BLN14, WL8);
sram_cell_6t_3 inst_cell_7_14 ( BL14, BLN14, WL7);
sram_cell_6t_3 inst_cell_6_14 ( BL14, BLN14, WL6);
sram_cell_6t_3 inst_cell_5_14 ( BL14, BLN14, WL5);
sram_cell_6t_3 inst_cell_4_14 ( BL14, BLN14, WL4);
sram_cell_6t_3 inst_cell_3_14 ( BL14, BLN14, WL3);
sram_cell_6t_3 inst_cell_2_14 ( BL14, BLN14, WL2);
sram_cell_6t_3 inst_cell_1_14 ( BL14, BLN14, WL1);
sram_cell_6t_3 inst_cell_0_14 ( BL14, BLN14, WL0);
sram_cell_6t_3 inst_cell_13_13 ( BL13, BLN13, WL13);
sram_cell_6t_3 inst_cell_12_13 ( BL13, BLN13, WL12);
sram_cell_6t_3 inst_cell_11_13 ( BL13, BLN13, WL11);
sram_cell_6t_3 inst_cell_10_13 ( BL13, BLN13, WL10);
sram_cell_6t_3 inst_cell_9_13 ( BL13, BLN13, WL9);
sram_cell_6t_3 inst_cell_8_13 ( BL13, BLN13, WL8);
sram_cell_6t_3 inst_cell_7_13 ( BL13, BLN13, WL7);
sram_cell_6t_3 inst_cell_6_13 ( BL13, BLN13, WL6);
sram_cell_6t_3 inst_cell_5_13 ( BL13, BLN13, WL5);
sram_cell_6t_3 inst_cell_4_13 ( BL13, BLN13, WL4);
sram_cell_6t_3 inst_cell_3_13 ( BL13, BLN13, WL3);
sram_cell_6t_3 inst_cell_2_13 ( BL13, BLN13, WL2);
sram_cell_6t_3 inst_cell_1_13 ( BL13, BLN13, WL1);
sram_cell_6t_3 inst_cell_0_13 ( BL13, BLN13, WL0);
sram_cell_6t_3 inst_cell_13_12 ( BL12, BLN12, WL13);
sram_cell_6t_3 inst_cell_12_12 ( BL12, BLN12, WL12);
sram_cell_6t_3 inst_cell_11_12 ( BL12, BLN12, WL11);
sram_cell_6t_3 inst_cell_10_12 ( BL12, BLN12, WL10);
sram_cell_6t_3 inst_cell_9_12 ( BL12, BLN12, WL9);
sram_cell_6t_3 inst_cell_8_12 ( BL12, BLN12, WL8);
sram_cell_6t_3 inst_cell_7_12 ( BL12, BLN12, WL7);
sram_cell_6t_3 inst_cell_6_12 ( BL12, BLN12, WL6);
sram_cell_6t_3 inst_cell_5_12 ( BL12, BLN12, WL5);
sram_cell_6t_3 inst_cell_4_12 ( BL12, BLN12, WL4);
sram_cell_6t_3 inst_cell_3_12 ( BL12, BLN12, WL3);
sram_cell_6t_3 inst_cell_2_12 ( BL12, BLN12, WL2);
sram_cell_6t_3 inst_cell_1_12 ( BL12, BLN12, WL1);
sram_cell_6t_3 inst_cell_0_12 ( BL12, BLN12, WL0);
sram_cell_6t_3 inst_cell_13_11 ( BL11, BLN11, WL13);
sram_cell_6t_3 inst_cell_12_11 ( BL11, BLN11, WL12);
sram_cell_6t_3 inst_cell_11_11 ( BL11, BLN11, WL11);
sram_cell_6t_3 inst_cell_10_11 ( BL11, BLN11, WL10);
sram_cell_6t_3 inst_cell_9_11 ( BL11, BLN11, WL9);
sram_cell_6t_3 inst_cell_8_11 ( BL11, BLN11, WL8);
sram_cell_6t_3 inst_cell_7_11 ( BL11, BLN11, WL7);
sram_cell_6t_3 inst_cell_6_11 ( BL11, BLN11, WL6);
sram_cell_6t_3 inst_cell_5_11 ( BL11, BLN11, WL5);
sram_cell_6t_3 inst_cell_4_11 ( BL11, BLN11, WL4);
sram_cell_6t_3 inst_cell_3_11 ( BL11, BLN11, WL3);
sram_cell_6t_3 inst_cell_2_11 ( BL11, BLN11, WL2);
sram_cell_6t_3 inst_cell_1_11 ( BL11, BLN11, WL1);
sram_cell_6t_3 inst_cell_0_11 ( BL11, BLN11, WL0);
sram_cell_6t_3 inst_cell_13_10 ( BL10, BLN10, WL13);
sram_cell_6t_3 inst_cell_12_10 ( BL10, BLN10, WL12);
sram_cell_6t_3 inst_cell_11_10 ( BL10, BLN10, WL11);
sram_cell_6t_3 inst_cell_10_10 ( BL10, BLN10, WL10);
sram_cell_6t_3 inst_cell_9_10 ( BL10, BLN10, WL9);
sram_cell_6t_3 inst_cell_8_10 ( BL10, BLN10, WL8);
sram_cell_6t_3 inst_cell_7_10 ( BL10, BLN10, WL7);
sram_cell_6t_3 inst_cell_6_10 ( BL10, BLN10, WL6);
sram_cell_6t_3 inst_cell_5_10 ( BL10, BLN10, WL5);
sram_cell_6t_3 inst_cell_4_10 ( BL10, BLN10, WL4);
sram_cell_6t_3 inst_cell_3_10 ( BL10, BLN10, WL3);
sram_cell_6t_3 inst_cell_2_10 ( BL10, BLN10, WL2);
sram_cell_6t_3 inst_cell_1_10 ( BL10, BLN10, WL1);
sram_cell_6t_3 inst_cell_0_10 ( BL10, BLN10, WL0);
sram_cell_6t_3 inst_cell_13_9 ( BL9, BLN9, WL13);
sram_cell_6t_3 inst_cell_12_9 ( BL9, BLN9, WL12);
sram_cell_6t_3 inst_cell_11_9 ( BL9, BLN9, WL11);
sram_cell_6t_3 inst_cell_10_9 ( BL9, BLN9, WL10);
sram_cell_6t_3 inst_cell_9_9 ( BL9, BLN9, WL9);
sram_cell_6t_3 inst_cell_8_9 ( BL9, BLN9, WL8);
sram_cell_6t_3 inst_cell_7_9 ( BL9, BLN9, WL7);
sram_cell_6t_3 inst_cell_6_9 ( BL9, BLN9, WL6);
sram_cell_6t_3 inst_cell_5_9 ( BL9, BLN9, WL5);
sram_cell_6t_3 inst_cell_4_9 ( BL9, BLN9, WL4);
sram_cell_6t_3 inst_cell_3_9 ( BL9, BLN9, WL3);
sram_cell_6t_3 inst_cell_2_9 ( BL9, BLN9, WL2);
sram_cell_6t_3 inst_cell_1_9 ( BL9, BLN9, WL1);
sram_cell_6t_3 inst_cell_0_9 ( BL9, BLN9, WL0);
sram_cell_6t_3 inst_cell_13_8 ( BL8, BLN8, WL13);
sram_cell_6t_3 inst_cell_12_8 ( BL8, BLN8, WL12);
sram_cell_6t_3 inst_cell_11_8 ( BL8, BLN8, WL11);
sram_cell_6t_3 inst_cell_10_8 ( BL8, BLN8, WL10);
sram_cell_6t_3 inst_cell_9_8 ( BL8, BLN8, WL9);
sram_cell_6t_3 inst_cell_8_8 ( BL8, BLN8, WL8);
sram_cell_6t_3 inst_cell_7_8 ( BL8, BLN8, WL7);
sram_cell_6t_3 inst_cell_6_8 ( BL8, BLN8, WL6);
sram_cell_6t_3 inst_cell_5_8 ( BL8, BLN8, WL5);
sram_cell_6t_3 inst_cell_4_8 ( BL8, BLN8, WL4);
sram_cell_6t_3 inst_cell_3_8 ( BL8, BLN8, WL3);
sram_cell_6t_3 inst_cell_2_8 ( BL8, BLN8, WL2);
sram_cell_6t_3 inst_cell_1_8 ( BL8, BLN8, WL1);
sram_cell_6t_3 inst_cell_0_8 ( BL8, BLN8, WL0);
sram_cell_6t_3 inst_cell_13_7 ( BL7, BLN7, WL13);
sram_cell_6t_3 inst_cell_12_7 ( BL7, BLN7, WL12);
sram_cell_6t_3 inst_cell_11_7 ( BL7, BLN7, WL11);
sram_cell_6t_3 inst_cell_10_7 ( BL7, BLN7, WL10);
sram_cell_6t_3 inst_cell_9_7 ( BL7, BLN7, WL9);
sram_cell_6t_3 inst_cell_8_7 ( BL7, BLN7, WL8);
sram_cell_6t_3 inst_cell_7_7 ( BL7, BLN7, WL7);
sram_cell_6t_3 inst_cell_6_7 ( BL7, BLN7, WL6);
sram_cell_6t_3 inst_cell_5_7 ( BL7, BLN7, WL5);
sram_cell_6t_3 inst_cell_4_7 ( BL7, BLN7, WL4);
sram_cell_6t_3 inst_cell_3_7 ( BL7, BLN7, WL3);
sram_cell_6t_3 inst_cell_2_7 ( BL7, BLN7, WL2);
sram_cell_6t_3 inst_cell_1_7 ( BL7, BLN7, WL1);
sram_cell_6t_3 inst_cell_0_7 ( BL7, BLN7, WL0);
sram_cell_6t_3 inst_cell_13_6 ( BL6, BLN6, WL13);
sram_cell_6t_3 inst_cell_12_6 ( BL6, BLN6, WL12);
sram_cell_6t_3 inst_cell_11_6 ( BL6, BLN6, WL11);
sram_cell_6t_3 inst_cell_10_6 ( BL6, BLN6, WL10);
sram_cell_6t_3 inst_cell_9_6 ( BL6, BLN6, WL9);
sram_cell_6t_3 inst_cell_8_6 ( BL6, BLN6, WL8);
sram_cell_6t_3 inst_cell_7_6 ( BL6, BLN6, WL7);
sram_cell_6t_3 inst_cell_6_6 ( BL6, BLN6, WL6);
sram_cell_6t_3 inst_cell_5_6 ( BL6, BLN6, WL5);
sram_cell_6t_3 inst_cell_4_6 ( BL6, BLN6, WL4);
sram_cell_6t_3 inst_cell_3_6 ( BL6, BLN6, WL3);
sram_cell_6t_3 inst_cell_2_6 ( BL6, BLN6, WL2);
sram_cell_6t_3 inst_cell_1_6 ( BL6, BLN6, WL1);
sram_cell_6t_3 inst_cell_0_6 ( BL6, BLN6, WL0);
sram_cell_6t_3 inst_cell_13_5 ( BL5, BLN5, WL13);
sram_cell_6t_3 inst_cell_12_5 ( BL5, BLN5, WL12);
sram_cell_6t_3 inst_cell_11_5 ( BL5, BLN5, WL11);
sram_cell_6t_3 inst_cell_10_5 ( BL5, BLN5, WL10);
sram_cell_6t_3 inst_cell_9_5 ( BL5, BLN5, WL9);
sram_cell_6t_3 inst_cell_8_5 ( BL5, BLN5, WL8);
sram_cell_6t_3 inst_cell_7_5 ( BL5, BLN5, WL7);
sram_cell_6t_3 inst_cell_6_5 ( BL5, BLN5, WL6);
sram_cell_6t_3 inst_cell_5_5 ( BL5, BLN5, WL5);
sram_cell_6t_3 inst_cell_4_5 ( BL5, BLN5, WL4);
sram_cell_6t_3 inst_cell_3_5 ( BL5, BLN5, WL3);
sram_cell_6t_3 inst_cell_2_5 ( BL5, BLN5, WL2);
sram_cell_6t_3 inst_cell_1_5 ( BL5, BLN5, WL1);
sram_cell_6t_3 inst_cell_0_5 ( BL5, BLN5, WL0);
sram_cell_6t_3 inst_cell_13_4 ( BL4, BLN4, WL13);
sram_cell_6t_3 inst_cell_12_4 ( BL4, BLN4, WL12);
sram_cell_6t_3 inst_cell_11_4 ( BL4, BLN4, WL11);
sram_cell_6t_3 inst_cell_10_4 ( BL4, BLN4, WL10);
sram_cell_6t_3 inst_cell_9_4 ( BL4, BLN4, WL9);
sram_cell_6t_3 inst_cell_8_4 ( BL4, BLN4, WL8);
sram_cell_6t_3 inst_cell_7_4 ( BL4, BLN4, WL7);
sram_cell_6t_3 inst_cell_6_4 ( BL4, BLN4, WL6);
sram_cell_6t_3 inst_cell_5_4 ( BL4, BLN4, WL5);
sram_cell_6t_3 inst_cell_4_4 ( BL4, BLN4, WL4);
sram_cell_6t_3 inst_cell_3_4 ( BL4, BLN4, WL3);
sram_cell_6t_3 inst_cell_2_4 ( BL4, BLN4, WL2);
sram_cell_6t_3 inst_cell_1_4 ( BL4, BLN4, WL1);
sram_cell_6t_3 inst_cell_0_4 ( BL4, BLN4, WL0);
sram_cell_6t_3 inst_cell_13_3 ( BL3, BLN3, WL13);
sram_cell_6t_3 inst_cell_12_3 ( BL3, BLN3, WL12);
sram_cell_6t_3 inst_cell_11_3 ( BL3, BLN3, WL11);
sram_cell_6t_3 inst_cell_10_3 ( BL3, BLN3, WL10);
sram_cell_6t_3 inst_cell_9_3 ( BL3, BLN3, WL9);
sram_cell_6t_3 inst_cell_8_3 ( BL3, BLN3, WL8);
sram_cell_6t_3 inst_cell_7_3 ( BL3, BLN3, WL7);
sram_cell_6t_3 inst_cell_6_3 ( BL3, BLN3, WL6);
sram_cell_6t_3 inst_cell_5_3 ( BL3, BLN3, WL5);
sram_cell_6t_3 inst_cell_4_3 ( BL3, BLN3, WL4);
sram_cell_6t_3 inst_cell_3_3 ( BL3, BLN3, WL3);
sram_cell_6t_3 inst_cell_2_3 ( BL3, BLN3, WL2);
sram_cell_6t_3 inst_cell_1_3 ( BL3, BLN3, WL1);
sram_cell_6t_3 inst_cell_0_3 ( BL3, BLN3, WL0);
sram_cell_6t_3 inst_cell_13_2 ( BL2, BLN2, WL13);
sram_cell_6t_3 inst_cell_12_2 ( BL2, BLN2, WL12);
sram_cell_6t_3 inst_cell_11_2 ( BL2, BLN2, WL11);
sram_cell_6t_3 inst_cell_10_2 ( BL2, BLN2, WL10);
sram_cell_6t_3 inst_cell_9_2 ( BL2, BLN2, WL9);
sram_cell_6t_3 inst_cell_8_2 ( BL2, BLN2, WL8);
sram_cell_6t_3 inst_cell_7_2 ( BL2, BLN2, WL7);
sram_cell_6t_3 inst_cell_6_2 ( BL2, BLN2, WL6);
sram_cell_6t_3 inst_cell_5_2 ( BL2, BLN2, WL5);
sram_cell_6t_3 inst_cell_4_2 ( BL2, BLN2, WL4);
sram_cell_6t_3 inst_cell_3_2 ( BL2, BLN2, WL3);
sram_cell_6t_3 inst_cell_2_2 ( BL2, BLN2, WL2);
sram_cell_6t_3 inst_cell_1_2 ( BL2, BLN2, WL1);
sram_cell_6t_3 inst_cell_0_2 ( BL2, BLN2, WL0);
sram_cell_6t_3 inst_cell_13_1 ( BL1, BLN1, WL13);
sram_cell_6t_3 inst_cell_13_0 ( BL0, BLN0, WL13);
sram_cell_6t_3 inst_cell_12_1 ( BL1, BLN1, WL12);
sram_cell_6t_3 inst_cell_12_0 ( BL0, BLN0, WL12);
sram_cell_6t_3 inst_cell_11_1 ( BL1, BLN1, WL11);
sram_cell_6t_3 inst_cell_11_0 ( BL0, BLN0, WL11);
sram_cell_6t_3 inst_cell_10_1 ( BL1, BLN1, WL10);
sram_cell_6t_3 inst_cell_10_0 ( BL0, BLN0, WL10);
sram_cell_6t_3 inst_cell_9_1 ( BL1, BLN1, WL9);
sram_cell_6t_3 inst_cell_9_0 ( BL0, BLN0, WL9);
sram_cell_6t_3 inst_cell_8_1 ( BL1, BLN1, WL8);
sram_cell_6t_3 inst_cell_8_0 ( BL0, BLN0, WL8);
sram_cell_6t_3 inst_cell_7_1 ( BL1, BLN1, WL7);
sram_cell_6t_3 inst_cell_7_0 ( BL0, BLN0, WL7);
sram_cell_6t_3 inst_cell_6_1 ( BL1, BLN1, WL6);
sram_cell_6t_3 inst_cell_6_0 ( BL0, BLN0, WL6);
sram_cell_6t_3 inst_cell_5_1 ( BL1, BLN1, WL5);
sram_cell_6t_3 inst_cell_5_0 ( BL0, BLN0, WL5);
sram_cell_6t_3 inst_cell_4_1 ( BL1, BLN1, WL4);
sram_cell_6t_3 inst_cell_4_0 ( BL0, BLN0, WL4);
sram_cell_6t_3 inst_cell_3_1 ( BL1, BLN1, WL3);
sram_cell_6t_3 inst_cell_3_0 ( BL0, BLN0, WL3);
sram_cell_6t_3 inst_cell_2_1 ( BL1, BLN1, WL2);
sram_cell_6t_3 inst_cell_2_0 ( BL0, BLN0, WL2);
sram_cell_6t_3 inst_cell_1_1 ( BL1, BLN1, WL1);
sram_cell_6t_3 inst_cell_0_1 ( BL1, BLN1, WL0);
sram_cell_6t_3 inst_cell_1_0 ( BL0, BLN0, WL1);
sram_cell_6t_3 inst_cell_0_0 ( BL0, BLN0, WL0);
sram_cell_6t_3 inst_cell_5_95 ( BL95, BLN95, WL5);
sram_cell_6t_3 inst_cell_4_95 ( BL95, BLN95, WL4);
sram_cell_6t_3 inst_cell_3_95 ( BL95, BLN95, WL3);
sram_cell_6t_3 inst_cell_2_95 ( BL95, BLN95, WL2);
sram_cell_6t_3 inst_cell_1_95 ( BL95, BLN95, WL1);
sram_cell_6t_3 inst_cell_0_95 ( BL95, BLN95, WL0);
sram_cell_6t_3 inst_cell_5_62 ( BL62, BLN62, WL5);
sram_cell_6t_3 inst_cell_5_29 ( BL29, BLN29, WL5);
sram_cell_6t_3 inst_cell_4_62 ( BL62, BLN62, WL4);
sram_cell_6t_3 inst_cell_4_29 ( BL29, BLN29, WL4);
sram_cell_6t_3 inst_cell_3_62 ( BL62, BLN62, WL3);
sram_cell_6t_3 inst_cell_3_29 ( BL29, BLN29, WL3);
sram_cell_6t_3 inst_cell_2_62 ( BL62, BLN62, WL2);
sram_cell_6t_3 inst_cell_2_29 ( BL29, BLN29, WL2);
sram_cell_6t_3 inst_cell_1_62 ( BL62, BLN62, WL1);
sram_cell_6t_3 inst_cell_0_62 ( BL62, BLN62, WL0);
sram_cell_6t_3 inst_cell_1_29 ( BL29, BLN29, WL1);
sram_cell_6t_3 inst_cell_0_29 ( BL29, BLN29, WL0);
inverter_compiler inst_invComp ( clk_bar, clk);
sense_amp_clocked_compiler inst_senAmp7 ( dout7, net21306, DL7, DLN7,
     sense_en);
sense_amp_clocked_compiler inst_senAmp6 ( dout6, net21307, DL6, DLN6,
     sense_en);
sense_amp_clocked_compiler inst_senAmp5 ( dout5, net21308, DL5, DLN5,
     sense_en);
sense_amp_clocked_compiler inst_senAmp4 ( dout4, net21309, DL4, DLN4,
     sense_en);
sense_amp_clocked_compiler inst_senAmp3 ( dout3, net21310, DL3, DLN3,
     sense_en);
sense_amp_clocked_compiler inst_senAmp2 ( dout2, net21311, DL2, DLN2,
     sense_en);
sense_amp_clocked_compiler inst_senAmp0 ( dout0, net21312, DL0, DLN0,
     sense_en);
sense_amp_clocked_compiler inst_senAmp1 ( dout1, net21313, DL1, DLN1,
     sense_en);
write_driver_compiler inst_writeDriver7 ( DL7, DLN7, clk_bar, din7,
     write_en);
write_driver_compiler inst_writeDriver6 ( DL6, DLN6, clk_bar, din6,
     write_en);
write_driver_compiler inst_writeDriver5 ( DL5, DLN5, clk_bar, din5,
     write_en);
write_driver_compiler inst_writeDriver4 ( DL4, DLN4, clk_bar, din4,
     write_en);
write_driver_compiler inst_writeDriver3 ( DL3, DLN3, clk_bar, din3,
     write_en);
write_driver_compiler inst_writeDriver2 ( DL2, DLN2, clk_bar, din2,
     write_en);
write_driver_compiler inst_writeDriver0 ( DL0, DLN0, clk_bar, din0,
     write_en);
write_driver_compiler inst_writeDriver1 ( DL1, DLN1, clk_bar, din1,
     write_en);
colDecoder inst_colDec ( .YF15(SL15), .YF14(SL14), .YF13(SL13),
     .YF12(SL12), .YF11(SL11), .YF10(SL10), .YF9(SL9), .YF8(SL8),
     .YF7(SL7), .YF6(SL6), .YF5(SL5), .YF4(SL4), .YF3(SL3), .YF2(SL2),
     .YF1(SL1), .YF0(SL0), .CLK(clk_bar), .A3_inv(inv_addr10),
     .A3(addr10), .A2_inv(inv_addr9), .A2(addr9), .A1_inv(inv_addr8),
     .A1(addr8), .A0_inv(inv_addr7), .A0(addr7));
invCol inst_invCol ( .Abar3(inv_addr10), .Abar2(inv_addr9),
     .Abar1(inv_addr8), .Abar0(inv_addr7), .A3(addr10), .A2(addr9),
     .A1(addr8), .A0(addr7));
precharge_compiler inst_precharge127 ( BL127, BLN127, clk_bar);
precharge_compiler inst_precharge126 ( BL126, BLN126, clk_bar);
precharge_compiler inst_precharge125 ( BL125, BLN125, clk_bar);
precharge_compiler inst_precharge124 ( BL124, BLN124, clk_bar);
precharge_compiler inst_precharge123 ( BL123, BLN123, clk_bar);
precharge_compiler inst_precharge122 ( BL122, BLN122, clk_bar);
precharge_compiler inst_precharge121 ( BL121, BLN121, clk_bar);
precharge_compiler inst_precharge120 ( BL120, BLN120, clk_bar);
precharge_compiler inst_precharge119 ( BL119, BLN119, clk_bar);
precharge_compiler inst_precharge118 ( BL118, BLN118, clk_bar);
precharge_compiler inst_precharge117 ( BL117, BLN117, clk_bar);
precharge_compiler inst_precharge116 ( BL116, BLN116, clk_bar);
precharge_compiler inst_precharge115 ( BL115, BLN115, clk_bar);
precharge_compiler inst_precharge114 ( BL114, BLN114, clk_bar);
precharge_compiler inst_precharge113 ( BL113, BLN113, clk_bar);
precharge_compiler inst_precharge112 ( BL112, BLN112, clk_bar);
precharge_compiler inst_precharge111 ( BL111, BLN111, clk_bar);
precharge_compiler inst_precharge110 ( BL110, BLN110, clk_bar);
precharge_compiler inst_precharge109 ( BL109, BLN109, clk_bar);
precharge_compiler inst_precharge108 ( BL108, BLN108, clk_bar);
precharge_compiler inst_precharge107 ( BL107, BLN107, clk_bar);
precharge_compiler inst_precharge106 ( BL106, BLN106, clk_bar);
precharge_compiler inst_precharge105 ( BL105, BLN105, clk_bar);
precharge_compiler inst_precharge104 ( BL104, BLN104, clk_bar);
precharge_compiler inst_precharge103 ( BL103, BLN103, clk_bar);
precharge_compiler inst_precharge102 ( BL102, BLN102, clk_bar);
precharge_compiler inst_precharge101 ( BL101, BLN101, clk_bar);
precharge_compiler inst_precharge100 ( BL100, BLN100, clk_bar);
precharge_compiler inst_precharge99 ( BL99, BLN99, clk_bar);
precharge_compiler inst_precharge98 ( BL98, BLN98, clk_bar);
precharge_compiler inst_precharge97 ( BL97, BLN97, clk_bar);
precharge_compiler inst_precharge96 ( BL96, BLN96, clk_bar);
precharge_compiler inst_precharge95 ( BL95, BLN95, clk_bar);
precharge_compiler inst_precharge94 ( BL94, BLN94, clk_bar);
precharge_compiler inst_precharge93 ( BL93, BLN93, clk_bar);
precharge_compiler inst_precharge92 ( BL92, BLN92, clk_bar);
precharge_compiler inst_precharge91 ( BL91, BLN91, clk_bar);
precharge_compiler inst_precharge90 ( BL90, BLN90, clk_bar);
precharge_compiler inst_precharge89 ( BL89, BLN89, clk_bar);
precharge_compiler inst_precharge88 ( BL88, BLN88, clk_bar);
precharge_compiler inst_precharge87 ( BL87, BLN87, clk_bar);
precharge_compiler inst_precharge86 ( BL86, BLN86, clk_bar);
precharge_compiler inst_precharge85 ( BL85, BLN85, clk_bar);
precharge_compiler inst_precharge84 ( BL84, BLN84, clk_bar);
precharge_compiler inst_precharge83 ( BL83, BLN83, clk_bar);
precharge_compiler inst_precharge82 ( BL82, BLN82, clk_bar);
precharge_compiler inst_precharge81 ( BL81, BLN81, clk_bar);
precharge_compiler inst_precharge80 ( BL80, BLN80, clk_bar);
precharge_compiler inst_precharge79 ( BL79, BLN79, clk_bar);
precharge_compiler inst_precharge78 ( BL78, BLN78, clk_bar);
precharge_compiler inst_precharge77 ( BL77, BLN77, clk_bar);
precharge_compiler inst_precharge76 ( BL76, BLN76, clk_bar);
precharge_compiler inst_precharge75 ( BL75, BLN75, clk_bar);
precharge_compiler inst_precharge74 ( BL74, BLN74, clk_bar);
precharge_compiler inst_precharge73 ( BL73, BLN73, clk_bar);
precharge_compiler inst_precharge72 ( BL72, BLN72, clk_bar);
precharge_compiler inst_precharge71 ( BL71, BLN71, clk_bar);
precharge_compiler inst_precharge70 ( BL70, BLN70, clk_bar);
precharge_compiler inst_precharge69 ( BL69, BLN69, clk_bar);
precharge_compiler inst_precharge68 ( BL68, BLN68, clk_bar);
precharge_compiler inst_precharge67 ( BL67, BLN67, clk_bar);
precharge_compiler inst_precharge66 ( BL66, BLN66, clk_bar);
precharge_compiler inst_precharge65 ( BL65, BLN65, clk_bar);
precharge_compiler inst_precharge64 ( BL64, BLN64, clk_bar);
precharge_compiler inst_precharge63 ( BL63, BLN63, clk_bar);
precharge_compiler inst_precharge62 ( BL62, BLN62, clk_bar);
precharge_compiler inst_precharge61 ( BL61, BLN61, clk_bar);
precharge_compiler inst_precharge60 ( BL60, BLN60, clk_bar);
precharge_compiler inst_precharge59 ( BL59, BLN59, clk_bar);
precharge_compiler inst_precharge58 ( BL58, BLN58, clk_bar);
precharge_compiler inst_precharge57 ( BL57, BLN57, clk_bar);
precharge_compiler inst_precharge56 ( BL56, BLN56, clk_bar);
precharge_compiler inst_precharge55 ( BL55, BLN55, clk_bar);
precharge_compiler inst_precharge54 ( BL54, BLN54, clk_bar);
precharge_compiler inst_precharge53 ( BL53, BLN53, clk_bar);
precharge_compiler inst_precharge52 ( BL52, BLN52, clk_bar);
precharge_compiler inst_precharge51 ( BL51, BLN51, clk_bar);
precharge_compiler inst_precharge50 ( BL50, BLN50, clk_bar);
precharge_compiler inst_precharge49 ( BL49, BLN49, clk_bar);
precharge_compiler inst_precharge48 ( BL48, BLN48, clk_bar);
precharge_compiler inst_precharge47 ( BL47, BLN47, clk_bar);
precharge_compiler inst_precharge46 ( BL46, BLN46, clk_bar);
precharge_compiler inst_precharge45 ( BL45, BLN45, clk_bar);
precharge_compiler inst_precharge44 ( BL44, BLN44, clk_bar);
precharge_compiler inst_precharge43 ( BL43, BLN43, clk_bar);
precharge_compiler inst_precharge42 ( BL42, BLN42, clk_bar);
precharge_compiler inst_precharge41 ( BL41, BLN41, clk_bar);
precharge_compiler inst_precharge40 ( BL40, BLN40, clk_bar);
precharge_compiler inst_precharge39 ( BL39, BLN39, clk_bar);
precharge_compiler inst_precharge38 ( BL38, BLN38, clk_bar);
precharge_compiler inst_precharge37 ( BL37, BLN37, clk_bar);
precharge_compiler inst_precharge36 ( BL36, BLN36, clk_bar);
precharge_compiler inst_precharge35 ( BL35, BLN35, clk_bar);
precharge_compiler inst_precharge34 ( BL34, BLN34, clk_bar);
precharge_compiler inst_precharge33 ( BL33, BLN33, clk_bar);
precharge_compiler inst_precharge32 ( BL32, BLN32, clk_bar);
precharge_compiler inst_precharge31 ( BL31, BLN31, clk_bar);
precharge_compiler inst_precharge30 ( BL30, BLN30, clk_bar);
precharge_compiler inst_precharge29 ( BL29, BLN29, clk_bar);
precharge_compiler inst_precharge28 ( BL28, BLN28, clk_bar);
precharge_compiler inst_precharge27 ( BL27, BLN27, clk_bar);
precharge_compiler inst_precharge26 ( BL26, BLN26, clk_bar);
precharge_compiler inst_precharge25 ( BL25, BLN25, clk_bar);
precharge_compiler inst_precharge24 ( BL24, BLN24, clk_bar);
precharge_compiler inst_precharge23 ( BL23, BLN23, clk_bar);
precharge_compiler inst_precharge22 ( BL22, BLN22, clk_bar);
precharge_compiler inst_precharge21 ( BL21, BLN21, clk_bar);
precharge_compiler inst_precharge20 ( BL20, BLN20, clk_bar);
precharge_compiler inst_precharge19 ( BL19, BLN19, clk_bar);
precharge_compiler inst_precharge18 ( BL18, BLN18, clk_bar);
precharge_compiler inst_precharge17 ( BL17, BLN17, clk_bar);
precharge_compiler inst_precharge16 ( BL16, BLN16, clk_bar);
precharge_compiler inst_precharge15 ( BL15, BLN15, clk_bar);
precharge_compiler inst_precharge14 ( BL14, BLN14, clk_bar);
precharge_compiler inst_precharge13 ( BL13, BLN13, clk_bar);
precharge_compiler inst_precharge12 ( BL12, BLN12, clk_bar);
precharge_compiler inst_precharge11 ( BL11, BLN11, clk_bar);
precharge_compiler inst_precharge10 ( BL10, BLN10, clk_bar);
precharge_compiler inst_precharge9 ( BL9, BLN9, clk_bar);
precharge_compiler inst_precharge8 ( BL8, BLN8, clk_bar);
precharge_compiler inst_precharge7 ( BL7, BLN7, clk_bar);
precharge_compiler inst_precharge6 ( BL6, BLN6, clk_bar);
precharge_compiler inst_precharge5 ( BL5, BLN5, clk_bar);
precharge_compiler inst_precharge4 ( BL4, BLN4, clk_bar);
precharge_compiler inst_precharge3 ( BL3, BLN3, clk_bar);
precharge_compiler inst_precharge2 ( BL2, BLN2, clk_bar);
precharge_compiler inst_precharge1 ( BL1, BLN1, clk_bar);
precharge_compiler inst_precharge0 ( BL0, BLN0, clk_bar);
columnMux inst_colMux7 ( .Ybar(DLN7), .Y(DL7), .sel15(SL15),
     .sel14(SL14), .sel13(SL13), .sel12(SL12), .sel11(SL11),
     .sel10(SL10), .sel9(SL9), .sel8(SL8), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar15(BLN127), .A15(BL127), .Abar14(BLN126),
     .A14(BL126), .Abar13(BLN125), .A13(BL125), .Abar12(BLN124),
     .A12(BL124), .Abar11(BLN123), .A11(BL123), .Abar10(BLN122),
     .A10(BL122), .Abar9(BLN121), .A9(BL121), .Abar8(BLN120),
     .A8(BL120), .Abar7(BLN119), .A7(BL119), .Abar6(BLN118),
     .A6(BL118), .Abar5(BLN117), .A5(BL117), .Abar4(BLN116),
     .A4(BL116), .Abar3(BLN115), .A3(BL115), .Abar2(BLN114),
     .A2(BL114), .Abar1(BLN113), .A1(BL113), .Abar0(BLN112),
     .A0(BL112));
columnMux inst_colMux6 ( .Ybar(DLN6), .Y(DL6), .sel15(SL15),
     .sel14(SL14), .sel13(SL13), .sel12(SL12), .sel11(SL11),
     .sel10(SL10), .sel9(SL9), .sel8(SL8), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar15(BLN111), .A15(BL111), .Abar14(BLN110),
     .A14(BL110), .Abar13(BLN109), .A13(BL109), .Abar12(BLN108),
     .A12(BL108), .Abar11(BLN107), .A11(BL107), .Abar10(BLN106),
     .A10(BL106), .Abar9(BLN105), .A9(BL105), .Abar8(BLN104),
     .A8(BL104), .Abar7(BLN103), .A7(BL103), .Abar6(BLN102),
     .A6(BL102), .Abar5(BLN101), .A5(BL101), .Abar4(BLN100),
     .A4(BL100), .Abar3(BLN99), .A3(BL99), .Abar2(BLN98), .A2(BL98),
     .Abar1(BLN97), .A1(BL97), .Abar0(BLN96), .A0(BL96));
columnMux inst_colMux5 ( .Ybar(DLN5), .Y(DL5), .sel15(SL15),
     .sel14(SL14), .sel13(SL13), .sel12(SL12), .sel11(SL11),
     .sel10(SL10), .sel9(SL9), .sel8(SL8), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar15(BLN95), .A15(BL95), .Abar14(BLN94),
     .A14(BL94), .Abar13(BLN93), .A13(BL93), .Abar12(BLN92),
     .A12(BL92), .Abar11(BLN91), .A11(BL91), .Abar10(BLN90),
     .A10(BL90), .Abar9(BLN89), .A9(BL89), .Abar8(BLN88), .A8(BL88),
     .Abar7(BLN87), .A7(BL87), .Abar6(BLN86), .A6(BL86), .Abar5(BLN85),
     .A5(BL85), .Abar4(BLN84), .A4(BL84), .Abar3(BLN83), .A3(BL83),
     .Abar2(BLN82), .A2(BL82), .Abar1(BLN81), .A1(BL81), .Abar0(BLN80),
     .A0(BL80));
columnMux inst_colMux4 ( .Ybar(DLN4), .Y(DL4), .sel15(SL15),
     .sel14(SL14), .sel13(SL13), .sel12(SL12), .sel11(SL11),
     .sel10(SL10), .sel9(SL9), .sel8(SL8), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar15(BLN79), .A15(BL79), .Abar14(BLN78),
     .A14(BL78), .Abar13(BLN77), .A13(BL77), .Abar12(BLN76),
     .A12(BL76), .Abar11(BLN75), .A11(BL75), .Abar10(BLN74),
     .A10(BL74), .Abar9(BLN73), .A9(BL73), .Abar8(BLN72), .A8(BL72),
     .Abar7(BLN71), .A7(BL71), .Abar6(BLN70), .A6(BL70), .Abar5(BLN69),
     .A5(BL69), .Abar4(BLN68), .A4(BL68), .Abar3(BLN67), .A3(BL67),
     .Abar2(BLN66), .A2(BL66), .Abar1(BLN65), .A1(BL65), .Abar0(BLN64),
     .A0(BL64));
columnMux inst_colMux3 ( .Ybar(DLN3), .Y(DL3), .sel15(SL15),
     .sel14(SL14), .sel13(SL13), .sel12(SL12), .sel11(SL11),
     .sel10(SL10), .sel9(SL9), .sel8(SL8), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar15(BLN63), .A15(BL63), .Abar14(BLN62),
     .A14(BL62), .Abar13(BLN61), .A13(BL61), .Abar12(BLN60),
     .A12(BL60), .Abar11(BLN59), .A11(BL59), .Abar10(BLN58),
     .A10(BL58), .Abar9(BLN57), .A9(BL57), .Abar8(BLN56), .A8(BL56),
     .Abar7(BLN55), .A7(BL55), .Abar6(BLN54), .A6(BL54), .Abar5(BLN53),
     .A5(BL53), .Abar4(BLN52), .A4(BL52), .Abar3(BLN51), .A3(BL51),
     .Abar2(BLN50), .A2(BL50), .Abar1(BLN49), .A1(BL49), .Abar0(BLN48),
     .A0(BL48));
columnMux inst_colMux2 ( .Ybar(DLN2), .Y(DL2), .sel15(SL15),
     .sel14(SL14), .sel13(SL13), .sel12(SL12), .sel11(SL11),
     .sel10(SL10), .sel9(SL9), .sel8(SL8), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar15(BLN47), .A15(BL47), .Abar14(BLN46),
     .A14(BL46), .Abar13(BLN45), .A13(BL45), .Abar12(BLN44),
     .A12(BL44), .Abar11(BLN43), .A11(BL43), .Abar10(BLN42),
     .A10(BL42), .Abar9(BLN41), .A9(BL41), .Abar8(BLN40), .A8(BL40),
     .Abar7(BLN39), .A7(BL39), .Abar6(BLN38), .A6(BL38), .Abar5(BLN37),
     .A5(BL37), .Abar4(BLN36), .A4(BL36), .Abar3(BLN35), .A3(BL35),
     .Abar2(BLN34), .A2(BL34), .Abar1(BLN33), .A1(BL33), .Abar0(BLN32),
     .A0(BL32));
columnMux inst_colMux1 ( .Ybar(DLN1), .Y(DL1), .sel15(SL15),
     .sel14(SL14), .sel13(SL13), .sel12(SL12), .sel11(SL11),
     .sel10(SL10), .sel9(SL9), .sel8(SL8), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar15(BLN31), .A15(BL31), .Abar14(BLN30),
     .A14(BL30), .Abar13(BLN29), .A13(BL29), .Abar12(BLN28),
     .A12(BL28), .Abar11(BLN27), .A11(BL27), .Abar10(BLN26),
     .A10(BL26), .Abar9(BLN25), .A9(BL25), .Abar8(BLN24), .A8(BL24),
     .Abar7(BLN23), .A7(BL23), .Abar6(BLN22), .A6(BL22), .Abar5(BLN21),
     .A5(BL21), .Abar4(BLN20), .A4(BL20), .Abar3(BLN19), .A3(BL19),
     .Abar2(BLN18), .A2(BL18), .Abar1(BLN17), .A1(BL17), .Abar0(BLN16),
     .A0(BL16));
columnMux inst_colMux0 ( .Ybar(DLN0), .Y(DL0), .sel15(SL15),
     .sel14(SL14), .sel13(SL13), .sel12(SL12), .sel11(SL11),
     .sel10(SL10), .sel9(SL9), .sel8(SL8), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar15(BLN15), .A15(BL15), .Abar14(BLN14),
     .A14(BL14), .Abar13(BLN13), .A13(BL13), .Abar12(BLN12),
     .A12(BL12), .Abar11(BLN11), .A11(BL11), .Abar10(BLN10),
     .A10(BL10), .Abar9(BLN9), .A9(BL9), .Abar8(BLN8), .A8(BL8),
     .Abar7(BLN7), .A7(BL7), .Abar6(BLN6), .A6(BL6), .Abar5(BLN5),
     .A5(BL5), .Abar4(BLN4), .A4(BL4), .Abar3(BLN3), .A3(BL3),
     .Abar2(BLN2), .A2(BL2), .Abar1(BLN1), .A1(BL1), .Abar0(BLN0),
     .A0(BL0));
invRow inst_invRow ( .Abar6(inv_addr6), .Abar5(inv_addr5),
     .Abar4(inv_addr4), .Abar3(inv_addr3), .Abar2(inv_addr2),
     .Abar1(inv_addr1), .Abar0(inv_addr0), .A6(addr6), .A5(addr5),
     .A4(addr4), .A3(addr3), .A2(addr2), .A1(addr1), .A0(addr0));
rowDecoder inst_rowDec ( .YF127(WL127), .YF126(WL126), .YF125(WL125),
     .YF124(WL124), .YF123(WL123), .YF122(WL122), .YF121(WL121),
     .YF120(WL120), .YF119(WL119), .YF118(WL118), .YF117(WL117),
     .YF116(WL116), .YF115(WL115), .YF114(WL114), .YF113(WL113),
     .YF112(WL112), .YF111(WL111), .YF110(WL110), .YF109(WL109),
     .YF108(WL108), .YF107(WL107), .YF106(WL106), .YF105(WL105),
     .YF104(WL104), .YF103(WL103), .YF102(WL102), .YF101(WL101),
     .YF100(WL100), .YF99(WL99), .YF98(WL98), .YF97(WL97), .YF96(WL96),
     .YF95(WL95), .YF94(WL94), .YF93(WL93), .YF92(WL92), .YF91(WL91),
     .YF90(WL90), .YF89(WL89), .YF88(WL88), .YF87(WL87), .YF86(WL86),
     .YF85(WL85), .YF84(WL84), .YF83(WL83), .YF82(WL82), .YF81(WL81),
     .YF80(WL80), .YF79(WL79), .YF78(WL78), .YF77(WL77), .YF76(WL76),
     .YF75(WL75), .YF74(WL74), .YF73(WL73), .YF72(WL72), .YF71(WL71),
     .YF70(WL70), .YF69(WL69), .YF68(WL68), .YF67(WL67), .YF66(WL66),
     .YF65(WL65), .YF64(WL64), .YF63(WL63), .YF62(WL62), .YF61(WL61),
     .YF60(WL60), .YF59(WL59), .YF58(WL58), .YF57(WL57), .YF56(WL56),
     .YF55(WL55), .YF54(WL54), .YF53(WL53), .YF52(WL52), .YF51(WL51),
     .YF50(WL50), .YF49(WL49), .YF48(WL48), .YF47(WL47), .YF46(WL46),
     .YF45(WL45), .YF44(WL44), .YF43(WL43), .YF42(WL42), .YF41(WL41),
     .YF40(WL40), .YF39(WL39), .YF38(WL38), .YF37(WL37), .YF36(WL36),
     .YF35(WL35), .YF34(WL34), .YF33(WL33), .YF32(WL32), .YF31(WL31),
     .YF30(WL30), .YF29(WL29), .YF28(WL28), .YF27(WL27), .YF26(WL26),
     .YF25(WL25), .YF24(WL24), .YF23(WL23), .YF22(WL22), .YF21(WL21),
     .YF20(WL20), .YF19(WL19), .YF18(WL18), .YF17(WL17), .YF16(WL16),
     .YF15(WL15), .YF14(WL14), .YF13(WL13), .YF12(WL12), .YF11(WL11),
     .YF10(WL10), .YF9(WL9), .YF8(WL8), .YF7(WL7), .YF6(WL6),
     .YF5(WL5), .YF4(WL4), .YF3(WL3), .YF2(WL2), .YF1(WL1), .YF0(WL0),
     .CLK(clk_bar), .A6_inv(inv_addr6), .A6(addr6), .A5_inv(inv_addr5),
     .A5(addr5), .A4_inv(inv_addr4), .A4(addr4), .A3_inv(inv_addr3),
     .A3(addr3), .A2_inv(inv_addr2), .A2(addr2), .A1_inv(inv_addr1),
     .A1(addr1), .A0_inv(inv_addr0), .A0(addr0));

endmodule


// End HDL models
